`timescale 1ns / 1ps

`include "defines_riscv.v"

module tb_miriscv_alu();

parameter TEST_VALUES     = 10000;
parameter TIME_OPERATION  = 100;


wire [5:0]               operator_i;
wire [31:0]              operand_a_i;
wire [31:0]              operand_b_i;

wire [31:0]              result_o;
wire                     comparison_result_o;

alu_riscv DUT
(
  .ALUOp  (operator_i),
  .A      (operand_a_i),
  .B      (operand_b_i),

  .Result (result_o),
  .Flag   (comparison_result_o)
);

integer     i, err_count = 0;
reg [8*9:1] operator_type;

wire [31:0] result_dump;
wire        comparison_result_dump;

reg [103:0] running_line;

 assign operator_i             = running_line[103:98];
 assign comparison_result_dump = running_line[97];
 assign operand_a_i            = running_line[95:64];
 assign operand_b_i            = running_line[63:32];
 assign result_dump            = running_line[31:0];

initial
  begin
    $display( "Start test: ");
    
    for ( i = 0; i < TEST_VALUES; i = i + 1 )
      begin
        running_line = line_dump[i*104+:103];
        #TIME_OPERATION;
        if( (result_dump != result_o) || (comparison_result_dump != comparison_result_o) ) begin
          $display("ERROR Operator: %s", operator_type, " operand_A: %h", operand_a_i, " operand_B: %h", operand_b_i, " result_o: %h", result_o, " result_dump: %h", result_dump, " comparison_result_o: %h", comparison_result_o, " comparison_result_dump: %h", comparison_result_dump);
          err_count = err_count + 1'b1;
        end        
      end

    $display("Number of errors: %d", err_count);
    
    $stop;
  end
  
always @(*) begin
 case(operator_i)
   `ALU_ADD  : operator_type = "ALU_ADD  ";
   `ALU_SUB  : operator_type = "ALU_SUB  ";
   `ALU_XOR  : operator_type = "ALU_XOR  ";
   `ALU_OR   : operator_type = "ALU_OR   ";
   `ALU_AND  : operator_type = "ALU_AND  ";
   `ALU_SRA  : operator_type = "ALU_SRA  ";
   `ALU_SRL  : operator_type = "ALU_SRL  ";
   `ALU_SLL  : operator_type = "ALU_SLL  ";
   `ALU_LTS  : operator_type = "ALU_LTS  ";
   `ALU_LTU  : operator_type = "ALU_LTU  ";
   `ALU_GES  : operator_type = "ALU_GES  ";
   `ALU_GEU  : operator_type = "ALU_GEU  ";
   `ALU_EQ   : operator_type = "ALU_EQ   ";
   `ALU_NE   : operator_type = "ALU_NE   ";
   `ALU_SLTS : operator_type = "ALU_SLTS ";
   `ALU_SLTU : operator_type = "ALU_SLTU ";
   default   : operator_type = "NOP      ";
 endcase
end
  
reg [104*10000:0] line_dump = {
104'h0012153524c0895e81d29e93a5,
104'h308484d609b1f0566300000000,
104'h9c06b97b0d46df998d0699190d,
104'hbcb2c284658937521200000000,
104'h3000f3e30106d7cd0d00000000,
104'hbc3b23f1761e8dcd3d00000000,
104'h9076d457ed462df78c30f9a061,
104'h9c7cfde9f9e33724c6603520c0,
104'h94e2f784c5d513d2aa00000000,
104'h5472aff7e5bbd2727700000000,
104'hb88932d61247ecdb8f00000000,
104'hbc793069f2e77696ce00000000,
104'h04f4007ae8e2ca4ec500000000,
104'h9c2e58495cde8e28bd0e08081c,
104'h5496ab582db2a7266500000000,
104'h94b1ef62630573870a00000000,
104'h9cc03b22801064212000202000,
104'h30557845aacecccc9d00000000,
104'h60cb203e968983b81300000000,
104'h6086bc380da9a7d65300000000,
104'h08359fdd6beaa62ad500000000,
104'h0481174a02d7563eae00000000,
104'h940effe91de7c572cf00000000,
104'h60118449230509650a00000000,
104'h34e5730aca9e314c3cffffffff,
104'h347968bdf2452e618a00000000,
104'h0820c4b341ec4b34d800000000,
104'h003c20f378c48a128900ab0601,
104'h5475c50deb5b0265b600000000,
104'h54634bf9c6571513ae00000000,
104'h34de7502bc150fdd2affffffff,
104'h2885d79a0bb897be7100000000,
104'h0042f2418527f2554f6ae496d4,
104'h669dcc603b1d06333a00000000,
104'h04bf23327e0aaa4b1500000000,
104'h9478d99bf16c9c4bd900000000,
104'h30312307622635fb4c00000000,
104'h944fa1559f47b9a18f00000000,
104'h667c6da9f8dbcd60b700000000,
104'hb8cfc4569fae7d945c00000000,
104'h60adcbc05b44de378900000000,
104'h28a4ae3249e8233ed000000000,
104'hb8ebfec0d7a8c7fc5100000000,
104'h304b212f96061d7f0c00000000,
104'h94e12ccec26457edc800000000,
104'h08bb825a771ef2ed3d00000001,
104'hbc090cdb12bf05007e00000000,
104'h9036e5816d1cd9e7392a3c6654,
104'h660fd28f1fe9ebf6d300000000,
104'h3442d92f85bc14887800000000,
104'h2c2dda595b248b4b4900000000,
104'h909ff2ae3f150caf2a8afe0115,
104'h9c2c156358c33f388600152000,
104'h04c71a0c8ece2ff29c00000000,
104'h907d3599fa937dbc26ee4825dc,
104'h0439961773d18bb4a300000000,
104'h9c9799a82fd9d292b391908023,
104'h66afd8565f22290d4400000000,
104'h947bf8fdf7e59b36cb00000000,
104'h66f3091ae62d28db5a00000000,
104'h5414cfc129f682e2ed00000000,
104'h08ed536cdab29fb66500000000,
104'hb8da8ae2b5efbe94df00000000,
104'h003cf119792231ff445f2318bd,
104'h2ce8740cd015090b2a00000000,
104'h2855f6adab076fcf0e00000000,
104'h946e5daddccd5ebc9a00000000,
104'h04fedf72fde1f102c300000000,
104'h302b0eed562779e94e00000000,
104'h94b3d976678531340a00000000,
104'h345b6fb9b69c0e8a3800000000,
104'h663cd18779dc2bc4b800000000,
104'h044a74bf9449c65d9300000000,
104'h34823f2c04acb7ca59ffffffff,
104'h546dcb69dba6fcde4d00000000,
104'h906cb0b7d9b6a4266dda1491b4,
104'h90bb45e276653b49cade7eabbc,
104'h345b172db64a93719500000000,
104'hb8a3071a4602749b0400000000,
104'h087bd261f73498076900000000,
104'h08da6ebab444018d8800000001,
104'hbc147cd9289690042d00000000,
104'h2ce3c530c7975c9c2e00000000,
104'h308477e4080e41451c00000000,
104'h2cfea7a6fd149e072900000000,
104'h288e37901c4335678600000000,
104'h90ed3408da9eb7c63d7383cee7,
104'h04334ea766b855c47000000000,
104'h04b9f504735d7199ba00000000,
104'h042f3ab35e7d4779fa00000000,
104'h666a8e05d58d24f61a00000000,
104'h60dcf000b91b87613700000000,
104'hb84b273796603921c000000000,
104'h9c13259f26db461ab613041a26,
104'h2c3e99837d6e5f0fdc00000000,
104'h00436157863c03ff787f6556fe,
104'h043f5a9b7eed8d80db00000000,
104'h28e7c3b6cf3ced2b7900000000,
104'h34fd28e4fab0bcee61ffffffff,
104'h080b940917d0f578a100000000,
104'h0043779186a8639650ebdb27d6,
104'h007a8c59f59ab488351540e22a,
104'h00949a8a2960b175c1f54bffea,
104'h28e2e574c5cc01b49800000000,
104'h3025b27b4bb98c427300000000,
104'h34f622e6ecc550168affffffff,
104'h542758d14ed44b80a800000000,
104'h94549efda9d0ca8ca100000000,
104'h2c070bb90ef33466e600000000,
104'hb8cfd6c09f152fb52a00000000,
104'h60155a1d2ac6b5f48d00000000,
104'h664f75ff9e9c6de63800000000,
104'h04bccfa8796464e3c800000000,
104'hbc652345ca09ff411300000000,
104'hbc35a0c96be3b7aec700000000,
104'h945b0bddb65d059dba00000000,
104'h666216abc45c8295b900000000,
104'h2c492fd392da269ab400000000,
104'h343fbb3b7fc333908600000000,
104'h547d6df5faf92794f200000000,
104'h2c19452132dece5ebd00000000,
104'h08424fcd84f249a4e400000000,
104'h666543cfca54a879a900000000,
104'h90d095a8a14765a98e97f0012f,
104'h34fd8b6afb85e51e0bffffffff,
104'h90f78290ef64c83dc9934aad26,
104'h301b60e536bab1487500000000,
104'h66c7e8568f35cdbf6b00000000,
104'h344465e788d73fb4ae00000000,
104'h004df3819b493e45929731c72d,
104'h601444df289684e02d00000000,
104'h0425b75f4be169b0c200000000,
104'h2c8f1cf61e06b3050d00000000,
104'h2c7679fdec0c039d1800000000,
104'h5468ae1bd1c3761c8600000000,
104'hb8a0c024419dbf643b00000000,
104'h906c44f9d829efe95345ab108b,
104'h94ab196256adac225b00000000,
104'hbcf166fae28273e20400000000,
104'h5439ac0373ec50b4d800000000,
104'h08093e4d12dc0344b800000000,
104'h549c811239f287b6e500000000,
104'h60d0c5dca115890f2b00000000,
104'h3440905d81641b85c800000000,
104'h5413b5552750d5f9a100000000,
104'h668f8c6e1f82223a0400000000,
104'h662c2d2358cb5c809600000000,
104'h660a6e93148919b41200000000,
104'h94cb227096d8ace2b100000000,
104'h302ac2d555f6c38eed00000000,
104'h04158b2b2b7ab11bf500000000,
104'h3456b403ad93c1222700000000,
104'h604249ff84d3a8e4a700000000,
104'h60f3d7a6e7dcef90b900000000,
104'h2ca4da56496de5bbdb00000000,
104'hb864ba0fc92883b15100000000,
104'h2cd0bc5ea11546dd2a00000000,
104'h9c7d2a45faa2e6204520220040,
104'hbc41a10583be75427c00000000,
104'h66b9461472ff4f3cfe00000000,
104'h54b455f268b7dfaa6f00000000,
104'h6643460d86782321f000000000,
104'h2c1c7197382076914000000000,
104'h34940976287b0da9f6ffffffff,
104'h2ce2bf1ac5602831c000000000,
104'h283a625f741cde713900000000,
104'h9cd86a6ab01e1c873c18080230,
104'h2c1521932a3124d36200000000,
104'h600aec3515f0b14ee100000000,
104'h660be29d17a18bee4300000000,
104'h0464b5e3c9c336048600000000,
104'h301297cb2560f69dc100000000,
104'h90c69da28dad67e25a6bfa40d7,
104'h6003d62707165b7b2c00000000,
104'h00060a5d0cb8ade671beb8437d,
104'h9c9de17c3b5b60e5b619606432,
104'h04fbdfc2f7cf14ce9e00000000,
104'h90ae78585c2ab8f75584c0af09,
104'hb8902a3a20d00b12a000000000,
104'h3039600972da3d8cb400000000,
104'h666e8af5dd86dcf00d00000000,
104'h0825b0994bbccc427900000000,
104'h60cf63da9efef064fd00000000,
104'h08bde0d27b47e2738f00000001,
104'h5481c39a0371c129e300000000,
104'hb80e92431d58f93db100000000,
104'h3422119f44ca9cbc9500000000,
104'hbcf01d34e0f6a178ed00000000,
104'h94297a15527c1e5bf800000000,
104'h9046dcb78da95fc452ef8373df,
104'h284219e784236afd4600000000,
104'hb8c63a928c48487d9000000000,
104'h080beac117352d616a00000001,
104'h90427b5784d55bbcaa9720eb2e,
104'h903e6f0f7cb05202608e3d0d1c,
104'h2c5d4a4dbac5a1608b00000000,
104'h94d31dfea692831e2500000000,
104'h0419058332d10504a200000000,
104'h2ca48f7c498a64b01400000000,
104'h089ec9c03d25f2034b00000001,
104'h60ae68305c2390754700000000,
104'hbc433e97869caf7a3900000000,
104'h2cda058ab46851e5d000000000,
104'h349622502c467c458cffffffff,
104'h6603e9b707b522406a00000000,
104'h340895f911746affe800000000,
104'hb8a5e79e4b39e4817300000000,
104'h3076295bec11fe052300000000,
104'h00520eefa464e165c9b6f0556d,
104'h2c9ca70439ef8372df00000000,
104'h2cea5814d43383656700000000,
104'hbc4ea0419d583125b000000000,
104'h044110398224d2bf4900000000,
104'h34ecb91ad91000b720ffffffff,
104'h548e054c1c49b16f9300000000,
104'h9471b461e3954b822a00000000,
104'h9ce471f8c8aed72e5da4512848,
104'h301d3f9d3a4226a98400000000,
104'h9c95a9a82b1c8d7f3914892829,
104'h94897f1c12a97f005200000000,
104'hbc2c848959e82b96d000000000,
104'h08b759ea6e4bf5299700000001,
104'h046d8b87db535277a600000000,
104'h2c5d85d3bb80797c0000000000,
104'h0487e44c0fb4e8d66900000000,
104'h308653620c2ca8195900000000,
104'hbc62fd49c567d735cf00000000,
104'hb84839e590a8e4d85100000000,
104'h2cb4f9a4693b83cd7700000000,
104'hb82523654aec3758d800000000,
104'h284ddd4d9be20e9ac400000000,
104'h945c78b1b8dbe6f2b700000000,
104'h9cc378ee86984d5a3080484a00,
104'h663bed53775ad6c7b500000000,
104'h306a15f5d40387870700000000,
104'h903b0b977674a1ade94faa3a9f,
104'h6645e28b8b00f25f0100000000,
104'h086d808bdbc076428000000000,
104'h04611d9fc2e2ecdac500000000,
104'hb89827fa30d7b2e4af00000000,
104'h30b302da6657fbb9af00000000,
104'h94f4d86ee97c41aff800000000,
104'hbc8376ac06f78576ef00000000,
104'hbc70ef37e1cab47c9500000000,
104'h9cf7723eee304e4d6030420c60,
104'hbcf29c5ee59420ea2800000000,
104'h2c322f7d6414b4372900000000,
104'hb8f0eeaee1bbbc527700000000,
104'h083715156e40aaf58100000001,
104'h346a9fb9d53437d56800000000,
104'h28786271f0d57800aa00000000,
104'h9c079fc30ff8dc48f1009c4001,
104'h66be9bbc7d472e958e00000000,
104'h30f161dce21e664d3c00000000,
104'h60d4b5e6a977ebb1ef00000000,
104'h66ade7d05bd7a23caf00000000,
104'h2c25029b4a5cd20db900000000,
104'hbc098e2d1309c8351300000000,
104'h5432dc416528c6275100000000,
104'h90db983ab7cc98109917002a2e,
104'h949d12083ab8ea3a7100000000,
104'h2c317c0762f2356ae400000000,
104'h601513dd2abeda447d00000000,
104'h282cee5f5972c3a3e500000000,
104'h3076de6bede4a800c900000000,
104'h00a0aecc4157c1d1aff8709df0,
104'h00eda71cdbe696e8cdd43e05a8,
104'h6638139f708326d40600000000,
104'h54d14820a25e983dbd00000000,
104'h28b555de6a6e3d47dc00000000,
104'hb8a86c5e50bd86f47b00000000,
104'h30929d5825bc3f847800000000,
104'h2c7b7b89f6ae23ce5c00000000,
104'h2c11cc9b233cb3ab7900000000,
104'h90644605c8ddd146bbb9974373,
104'h90870cee0eb98794733e8b7a7d,
104'h040671030ce70f98ce00000000,
104'h286a1a61d4acecdc5900000000,
104'hbc5ca26fb9d9b8c0b300000000,
104'h9c7a4fbff4baf4e2753a44a274,
104'h66066cf10c9cfc7a3900000000,
104'h28017293028aecbe1500000000,
104'h6002fbf905271c434e00000000,
104'h00013f29025c7951b85db87aba,
104'h94847fb20846e7538d00000000,
104'h94d7b48eaf747331e800000000,
104'h28485909907af6abf500000000,
104'h28a620904c3d82bd7b00000000,
104'h04a005a64012a9032500000000,
104'h3486ebb60db87c1070ffffffff,
104'h5416cbf92d94ded82900000000,
104'h665e2551bc987b083000000000,
104'hbc60272dc02876695000000000,
104'hb8d0cf6aa126bf3f4d00000000,
104'hbcfaf32ef57a87aff500000000,
104'h60aeeacc5dca48129400000000,
104'h54b558a66a5e6065bc00000000,
104'h2cdc4308b8cf309c9e00000000,
104'h04fd7906fa23400b4600000000,
104'h2883fa6407c9cbbc9300000000,
104'h94aada74555bd3dbb700000000,
104'h6622d5f145b1800a6300000000,
104'h9cac93e0599372ce268012c000,
104'h00b44976688f63e41e43ad5a86,
104'h66c838f4902d19a55a00000000,
104'h040e43851c5c9967b900000000,
104'h6055861fab6826d9d000000000,
104'h0037b9656f6c6a6dd8a423d347,
104'h66a2cc884546d6a78d00000000,
104'h0445f3238b7e2491fc00000000,
104'h9c6e1e1fdcd27f0aa4421e0a84,
104'h040c978d1952b533a500000000,
104'h949f398e3ef98bc0f300000000,
104'h04ac782c5862056bc400000000,
104'h942e36435c033a450600000000,
104'h34cd1d509a0c161918ffffffff,
104'hbce2f066c55515d1aa00000000,
104'hbc0d12031a61dbd5c300000000,
104'h085934e9b20633630c00000000,
104'hb8f4f00ee961dafdc300000000,
104'h2c75ad73eb7c2db9f800000000,
104'h30792c03f24483ad8900000000,
104'h08378c736f0de14b1b00000000,
104'h00d6a128ad344dc1680aeeea15,
104'hb892f9122567e857cf00000000,
104'h0855dd8dab8d94d21b00000000,
104'h60c03b3e802ed6d95d00000000,
104'h2c412dfd828234420400000000,
104'h282ba7a5571b368b3600000000,
104'hbc196a0332bce3287900000000,
104'h9cf24baee48b42ec168242ac04,
104'h60d57fecaa605065c000000000,
104'h549759882e4665378c00000000,
104'h34b8c0c2717dfe8ffbffffffff,
104'hb85e5421bcee7068dc00000000,
104'h540bec5717e0e004c100000000,
104'h9075fb21eb5a9d3bb52f661a5e,
104'h60c4fd2e89c7b2e28f00000000,
104'h30dff6f6bfd8462ab000000000,
104'h90e9b49ad3eb1d02d602a99805,
104'h54c144cc820d63751a00000000,
104'h3038e6a771eb8804d700000000,
104'h5487628e0ef8c714f100000000,
104'hbc66861dcd02bd430500000000,
104'h340e3aeb1c4c18c79800000000,
104'h9cf67088ec9541d62a94408028,
104'h00b2d14a651b920537ce634f9c,
104'h2881fa3603ff729efe00000000,
104'h66feaddcfd9f7a0e3e00000000,
104'h28f43a34e8ba60387400000000,
104'h28580989b08361dc0600000000,
104'h3409164d12b46afc6800000000,
104'h60e2ba00c5ff202efe00000000,
104'h941b0f0d36799f09f300000000,
104'h047dddabfbb58d7c6b00000000,
104'hb80bcbbf1787d0360f00000000,
104'h948a47b6141500052a00000000,
104'h9cd3666ea6ea7626d4c2662684,
104'h94e5ac10cbb587c26b00000000,
104'h080277eb04fa4832f400000000,
104'h04468b618df0ea70e100000000,
104'h9c42e3bd85dc9974b940813481,
104'h94e4df16c9b05f8e6000000000,
104'h04a36432461e74cb3c00000000,
104'h9c1b855f372c0c555808045510,
104'h9c39d657738778d20e01505202,
104'h2c6e6d23dc183fc33000000000,
104'h606845f5d00073e50000000000,
104'h6621820f437c6e91f800000000,
104'h54d0b99aa129c01f5300000000,
104'h664c588f982fef3d5f00000000,
104'h90c3be9287fd5f5afa3ee1c87d,
104'h001699d12db8760270cf0fd39d,
104'h90b5b4e86b98d738312d63d05a,
104'h90892fc0120650df0c8f7f1f1e,
104'h0806db6b0d0acd131500000001,
104'h2c203107404a638d9400000000,
104'h342a1ba354c062028000000000,
104'h08098d1513e1e386c300000000,
104'hbcf695deedee4ee6dc00000000,
104'h54bc78107813d40d2700000000,
104'h08afed265f11c05b2300000001,
104'hbc5596ebab1c42173800000000,
104'h0011534d2264f2bdc976460aeb,
104'h2ce3eb4cc7c140628200000000,
104'h666754d7cee38e22c700000000,
104'hb8927fa4246da36fdb00000000,
104'hbc846514083ac26f7500000000,
104'h305ad31db58d7d721a00000000,
104'h2c1c2a1338c1233a8200000000,
104'h28ac05a058a85a6a5000000000,
104'h00d1889aa35243e3a423cc7e47,
104'h6032c3df65753c17ea00000000,
104'h0803703906aa13805400000000,
104'h66adf3405be455f0c800000000,
104'h90246739489bf8f237bf9fcb7f,
104'h047c1df3f8da8932b500000000,
104'h0828d6a95141aed58300000001,
104'h304d9ee39b1aa0dd3500000000,
104'h30581653b0fddf82fb00000000,
104'h34278dbb4f984da63000000000,
104'h9c8c38c418ee8118dd8c000018,
104'h04a36ae84630e20f6100000000,
104'h60ac9748592af1735500000000,
104'h66178b972f85ce500b00000000,
104'h9cef1deadee9d22cd3e91028d2,
104'h001445b12874dc69e989221b11,
104'h342c5779586aa4a1d500000000,
104'h9461dbe5c36a2c13d400000000,
104'h2852397da43f25ef7e00000000,
104'hb86b299dd687eec80f00000000,
104'h54c1b04483506aefa000000000,
104'h08c10f04825fe3cbbf00000001,
104'h5422eadb45bbbc3e7700000000,
104'h94229d0b45ba94107500000000,
104'h2cfc670af863323bc600000000,
104'h543601596ca84e585000000000,
104'h3018bd6331ce10fe9c00000000,
104'h04de325cbcd7e31eaf00000000,
104'hbc872d2c0eb4e4666900000000,
104'h08d95b40b2ef209ede00000001,
104'h2cc2e87485555c0faa00000000,
104'h281407f128610ed5c200000000,
104'h904d20099a69e751d324c75849,
104'h34dd111abafdeb7cfbffffffff,
104'h60c5cf728b61114dc200000000,
104'h54e64828cc38e6137100000000,
104'h944f49019e309cdb6100000000,
104'h2cbde3487bdf9bd0bf00000000,
104'h34c881bc91e06098c0ffffffff,
104'hbc2ca96359bf53b47e00000000,
104'h942a1d7354a8e2e25100000000,
104'h04a4de284973fa7de700000000,
104'hb8123aaf2441b5d58300000000,
104'h9cadee005b5cdea1b90cce0019,
104'h604afebf95bb934a7700000000,
104'h54f8da1af1732c5fe600000000,
104'h00d7e1aeaf0238e104da1a8fb3,
104'h28896460127e29b3fc00000000,
104'hb8d5ba48abe203f0c400000000,
104'h301ffb813fe13256c200000000,
104'hb8398a19732d4d9b5a00000000,
104'h66d066e4a0ff73cafe00000000,
104'hbc3a096b745d86b7bb00000000,
104'hbc7132bbe2f16948e200000000,
104'h60eff34cdfcc13e29800000000,
104'h044fdbed9f0817cb1000000000,
104'h34791189f25ee97bbd00000000,
104'h5455bc27ab5a0a0fb400000000,
104'h2caa08ac5444e79b8900000000,
104'h3089b5d413560c91ac00000000,
104'h2c1ae403351df61f3b00000000,
104'h949aa0243517a98d2f00000000,
104'h001a619934aae0a255c5423b89,
104'h9cde7302bcf964fef2d86002b0,
104'hb8d3fe36a7e0f280c100000000,
104'h00f23316e4a0b8a24192ebb925,
104'h54b4c16c69fd52d8fa00000000,
104'h9ce69dd0cd7fcff3ff668dd0cd,
104'h28dac986b5f42082e800000000,
104'h90a5955c4b89042e122c917259,
104'h901b978f37574e1dae4cd99299,
104'hb8fc4ca4f890184e2000000000,
104'h54ed1b50da913e022200000000,
104'h30763355ec9535122a00000000,
104'h9c3d7f5b7a0f1e511e0d1e511a,
104'hb8f4a1dae9f5a4f2eb00000000,
104'h0405b4f70bb704e26e00000000,
104'h08af455e5e3e502d7c00000001,
104'h2822c03145c5cb548b00000000,
104'h04094bd3121bf8bd3700000000,
104'h00c1c3d683f0ab00e1b26ed764,
104'hb8674fdfcea5365c4a00000000,
104'h006acd73d5669907cdd1667ba2,
104'h28f204eee4fa328cf400000000,
104'h04766153ec0d623f1a00000000,
104'h08f1a32ee3f62484ec00000001,
104'h9c79c681f31687472d10860121,
104'h042e138d5c6e8d45dd00000000,
104'h66f612c8ecc7d87a8f00000000,
104'h947fdbb3ff3c33857800000000,
104'h0055f6b9ab13d1f72769c8b0d2,
104'h007dca0ffb09dfc31387a9d30e,
104'h3006499b0c5db797bb00000000,
104'h9cf361cae6a4d83a49a0400a40,
104'hbc35557b6a8570f60a00000000,
104'h668c06d2184b1ce99600000000,
104'h2884e326091725712e00000000,
104'h66dee9d4bd3363896600000000,
104'h08bb0628763a98257500000001,
104'h66c7b43a8f4ad3959500000000,
104'h543da8cd7bbe43ea7c00000000,
104'h9cb7f4306fe4824cc9a4800049,
104'h2ce4d820c95a3761b400000000,
104'h9c6d48a5dad6aea8ad4408a088,
104'h946fcff1df06b0e30d00000000,
104'h30384d417041bd678300000000,
104'h00a8c6c451027a8d04ab415155,
104'hb8c0467280fcf504f900000000,
104'h540379ed06e5063aca00000000,
104'h66ef8d64df64f9bbc900000000,
104'h0042797584d84988b01ac2fe34,
104'h6674bc03e90809851000000000,
104'h666f3425ded659d0ac00000000,
104'h340498fb096bf823d700000000,
104'hb830c38f6186c8320d00000000,
104'h5448c3b791e9eb0ed300000000,
104'h084d77f99a17bd872f00000000,
104'h302720634e5bd583b700000000,
104'h90e32472c62ed66b5dcdf2199b,
104'h34ce03ec9c17b47f2fffffffff,
104'h30a22ac644cdbf3a9b00000000,
104'h34b1200062748abbe9ffffffff,
104'h901747832ec690128dd1d791a3,
104'h90632f07c6d51cb4aab633b36c,
104'h2cd01df0a01be8cf3700000000,
104'h66f8602ef0f46ca8e800000000,
104'h34e6841ccd68cd09d1ffffffff,
104'h305d8363bbeff692df00000000,
104'h603e8ed57d2c40215800000000,
104'h66cff5509f4bac2f9700000000,
104'h54835da20694a12e2900000000,
104'h00624b63c4ebb0f6d74dfc5a9b,
104'h08aea6d45d26c7134d00000001,
104'hb839bfc773bfd62a7f00000000,
104'h66a703744e5cdc65b900000000,
104'h66f05d64e09cd6c23900000000,
104'h2c40fb4f8118fb833100000000,
104'h0447ebef8f7f537dfe00000000,
104'h30aed0f05d878a880f00000000,
104'hb8199bcb33348ed56900000000,
104'h542b0da556cd57529a00000000,
104'h942e72295c24e9074900000000,
104'h9c69cd77d39d737a3a09417212,
104'h666c74f5d8bc1c0e7800000000,
104'h301ccb353992d0602500000000,
104'h288496d609ab37a85600000000,
104'h66962c682ce99b1cd300000000,
104'h040d633f1a005d510000000000,
104'h30560d5facf4588ee800000000,
104'h60b66a586cd03c40a000000000,
104'h600ecd251d68c14fd100000000,
104'h00006d0f00ed4d78daedba87da,
104'h006c1987d8605dbbc0cc774398,
104'h08a6490c4ce8cfb0d100000001,
104'h30a8bb0c51a8e1ee5100000000,
104'h94a2a4be45598367b300000000,
104'h94bf21067ec049c68000000000,
104'h607e5b53fc2426d74800000000,
104'h30c0ad808198b4dc3100000000,
104'h0453a8b5a741b1fd8300000000,
104'h349fc1423f00029100ffffffff,
104'h08b2158c643f52937e00000001,
104'h547887dff1472dfb8e00000000,
104'h944f234d9e742819e800000000,
104'h3024839b498569fa0a00000000,
104'h282fb81b5fa8bfc85100000000,
104'h9ca4d9864992fd282580d90001,
104'h94b64ae66cac509c5800000000,
104'h00af5d6c5e97dde22f473b4e8d,
104'h9cc1cf5a8313b7532701875203,
104'hbc6a5ddbd4ca0e449400000000,
104'h04c961e4921e32673c00000000,
104'h6023301b46b7b82a6f00000000,
104'h30a0b3ae417bde15f700000000,
104'hbc8b7c381639092f7200000000,
104'hbc5136a5a271f059e300000000,
104'h34c9490292e5ceb0cbffffffff,
104'h283409756898b4ee3100000000,
104'h6065c803cbaad1c85500000000,
104'h9c38a389712f49535e28010150,
104'hbce6e186cddaf356b500000000,
104'h0804410d08c118be8200000000,
104'h549f80983fd807f2b000000000,
104'h34560eefac9918303200000000,
104'h00029f05052f73fb5e32130063,
104'h90dc16d8b83ec2677de2d4bfc5,
104'hbc8511580ac6878a8d00000000,
104'h0464eb39c9f8d3d8f100000000,
104'h66da12deb4729a7fe500000000,
104'h041a13393411c6c52300000000,
104'h301691a32d18e8713100000000,
104'h282f36c55e5a0f27b400000000,
104'h66073a730e322cc16400000000,
104'h30320a8b642416b94800000000,
104'h34c544d88a4dfe879bffffffff,
104'h9ce6fbf4cdb5f8fa6ba4f8f049,
104'h0455ff23abf1eca2e300000000,
104'h545e9d2fbdecff24d900000000,
104'hbce11a58c2f059ace000000000,
104'h60afd1265f8edc361d00000000,
104'h90c9b64c9313180326daae4fb5,
104'h6682b7860584a8e80900000000,
104'h08b62d846cb5c5c06b00000000,
104'h085858bdb0fb9fb8f700000000,
104'h0852a151a5abe8c05700000000,
104'h603b11f3762798e34f00000000,
104'h605a45bdb48ecaa21d00000000,
104'h0043c1158723466346670778cd,
104'h54336d93664f14c19e00000000,
104'h541fb0d13f2a2ff55400000000,
104'h082a565f54a62c344c00000000,
104'hbc83449006286f135000000000,
104'h0416b46d2dc34ddc8600000000,
104'hbc3564836a5c2afdb800000000,
104'h28f7fecaef506a57a000000000,
104'h281fa98f3f84d4aa0900000000,
104'h90d47b42a8aac1fa557ebab8fd,
104'h088f49661edc22dcb800000001,
104'h28e70a62ceeb40e6d600000000,
104'hbc92c27025d4ce0aa900000000,
104'h00e7b374cf1a9af535024e6a04,
104'h662047dd405b0c73b600000000,
104'h30faf084f5ad27c45a00000000,
104'hbc70ed97e112ce112500000000,
104'h0893ba6027227eb14400000001,
104'h66bc944679cfb89e9f00000000,
104'h9c545493a864d2d3c944509388,
104'h9442955d8542e39d8500000000,
104'h54b9d96873440f098800000000,
104'h664b2f05969a54423400000000,
104'h661e85ed3d28b1f15100000000,
104'h088db0281b8e39901c00000001,
104'h085ec5ebbdda69e2b400000000,
104'h602764754e17e83f2f00000000,
104'h342cfff159f670fcec00000000,
104'h540f40551ece96ca9d00000000,
104'h66e02148c071a919e300000000,
104'h54b24cf664a5d9704b00000000,
104'h6648e9ff914277d78400000000,
104'hb824d4474989de2c1300000000,
104'h00d9f8e0b30e62911ce85b71cf,
104'h60144ced281568bb2a00000000,
104'h902e97795d776a61ee59fd18b3,
104'h6066065bcc5d8e95bb00000000,
104'h54bc461478652825ca00000000,
104'h302e94b75d8f32fa1e00000000,
104'hb83b07bd7665a879cb00000000,
104'h2c6dfcf1dbda42e4b400000000,
104'h34106e43200207bb0400000000,
104'h28bca0b279e6b110cd00000000,
104'hbcc9662c92a2ce004500000000,
104'h90d4ea6aa9cf31fc9e1bdb9637,
104'h086ec2cbdd600b2dc000000000,
104'h66a5b9424b5db7e1bb00000000,
104'h28408a2981d932d8b200000000,
104'hb8598d27b305aeb90b00000000,
104'h9424011148f0b860e100000000,
104'h607e72c5fcd7f844af00000000,
104'h08d0770ea0076adf0e00000001,
104'hb83aaf87756ca7ffd900000000,
104'h6686d26e0d1391312700000000,
104'h943a2d99747e7f21fc00000000,
104'h60dfdc3ebfafc5f25f00000000,
104'h34c0a7e881b428aa68ffffffff,
104'h30fd4c48fafd9380fb00000000,
104'h300c962119d33554a600000000,
104'h5429951b53f7cff6ef00000000,
104'h54f6d8aeed58d79db100000000,
104'h94b26ffe6490b9302100000000,
104'h087b24bdf6345fbf6800000000,
104'h348a290014b7d0ca6fffffffff,
104'h2c9530362a1f77b73e00000000,
104'h54fbaaeef723781f4600000000,
104'hbc9e9dca3dd01f40a000000000,
104'h947d4b53fa7a4c4df400000000,
104'h0019a8e3330067d7001a10ba33,
104'h006e567bdc38422d70a698a94c,
104'h049491aa2907f0b90f00000000,
104'h084b5b71966b825dd700000001,
104'h3011c911238322de0600000000,
104'h60a538004a2505394a00000000,
104'h9420dcbf41442d078800000000,
104'h9ce6e4b8cd38eedd7120e49841,
104'hbc9423222889bfac1300000000,
104'h2cb600e26caaab245500000000,
104'h947f2767fe37890d6f00000000,
104'h047a1e8bf4e0c9acc100000000,
104'h34e9d576d38c712218ffffffff,
104'h6056ce7fad7c99cff900000000,
104'h28646601c89295aa2500000000,
104'h60a46c48487186abe300000000,
104'h2c680a6fd04506218a00000000,
104'h90b3aa3667b83318700b992e17,
104'h083058ef60273fbf4e00000000,
104'hb867dd53cfb955b67200000000,
104'h90797869f2ca698294b311eb66,
104'h00f40968e84c54e198405e4a80,
104'h904f0c8f9e7c502bf8335ca466,
104'h66c6ad048de5a2b2cb00000000,
104'h28d7e1c6af1c222f3800000000,
104'h90704d75e050d909a120947c41,
104'h9cca594094d0ebcca1c0494080,
104'h0010c2c52112957f2523584446,
104'h66f594e6eb1dd3013b00000000,
104'h669743be2e4e156f9c00000000,
104'h600b6367169013842000000000,
104'h30e131eec2ca91f89500000000,
104'h6696ec2a2d02bad90500000000,
104'h5483a5a007745bf5e800000000,
104'h90cc1b609834243768f83f57f0,
104'h54cbb9e29775b801eb00000000,
104'h949bcdf2372934995200000000,
104'h3041987f83c37a788600000000,
104'h0438bd8d719a56bc3400000000,
104'hbcba460274b963787200000000,
104'h54f92c9af266371fcc00000000,
104'h9cc42db888223add4400289800,
104'hb841524b82c63ffa8c00000000,
104'h34fa6daef4c7ac408fffffffff,
104'h00e28688c5c0d54c81a35bd546,
104'h9c8ae2ac1565e2ffcb00e2ac01,
104'h941b2dfd361550d12a00000000,
104'h00faf442f59ee6363d99da7932,
104'h54236617469dbe003b00000000,
104'hbcf720bcee49b4c19300000000,
104'h90f27102e4e2561cc410271e20,
104'hbcb949247239213b7200000000,
104'h60a8e1aa515abc1db500000000,
104'h6651bd47a3566e01ac00000000,
104'h30cb87ba9798f8c03100000000,
104'h66df07b0beaba92e5700000000,
104'h603b1ba1765a3681b400000000,
104'h088079ac00b9c8a07300000001,
104'h0894aa8429393d9b7200000001,
104'h088f77461e3685f36d00000001,
104'h0066c259cd7eb00bfde57265ca,
104'h546b834dd70dfa7f1b00000000,
104'h28675dc5ce4b058b9600000000,
104'h54e50b48ca43fb658700000000,
104'h009690342d16479b2cacd7cf59,
104'h0812f3892511357d2200000000,
104'h04f9f1d4f3418d738300000000,
104'h601ee3173d580965b000000000,
104'h2c5ccb93b93638136c00000000,
104'h08544fbfa84d27799a00000000,
104'h90410319824eee339d0fed2a1f,
104'h307e4a0ffcefebd4df00000000,
104'hb8ecc6d4d98658500c00000000,
104'hbc600951c0ae7a545c00000000,
104'h0440f9f181a79ca84f00000000,
104'h9cd43790a8519a95a3501290a0,
104'h94c46058887c9b37f900000000,
104'h34defd9cbd0c53ef18ffffffff,
104'h040f8abb1f35e9b76b00000000,
104'h2cbecefe7d4b49839600000000,
104'h288582800b088fa31100000000,
104'h9cc7f6028f9fd6283f87d6000f,
104'h540535d70abd823a7b00000000,
104'h9496dfb62de2e87ec500000000,
104'h60ffa3aaffaee0765d00000000,
104'h60e527e6ca6b9ee1d700000000,
104'hbc1ec7a73d6eef15dd00000000,
104'h300d651b1af5a36aeb00000000,
104'h66694639d214d4932900000000,
104'h6009b4a3139347f82600000000,
104'h288ed88a1deb1528d600000000,
104'h6679068bf2c762268e00000000,
104'h08c9788892fbced2f700000001,
104'h66f7299aeea2e74e4500000000,
104'h047f4ce1feb6b5506d00000000,
104'h34d39764a782489004ffffffff,
104'h909154fc22acce1c593d9ae07b,
104'h90f3002ee6c68ec48d358eea6b,
104'h2c02d509051dec713b00000000,
104'h00679709cfa636884c0dcd921b,
104'h666581f3cbd3ed4ca700000000,
104'h300c1dbd18f1cc38e300000000,
104'hbc366d676c87b3680f00000000,
104'h902db0d95b6847f1d045f7288b,
104'h0017b1cd2fcbe34297e3950fc6,
104'hbc1053a720f7298cee00000000,
104'h0092de5425395f1772cc3d6b97,
104'hbcda3c32b40254a70400000000,
104'h94d022e8a05982e1b300000000,
104'h6031df4b638fac9e1f00000000,
104'h666e3c37dc8a205c1400000000,
104'h669abc7835f2708ce400000000,
104'h28671fa9ced73b04ae00000000,
104'h2c5cea0bb9525751a400000000,
104'h90ad676c5a8684180d2be37457,
104'h0483610a062a6b835400000000,
104'hbcee7e6adcd09690a100000000,
104'h603d09457a9ba7803700000000,
104'h08a58c544b03f32b0700000001,
104'h08ac8546592f51675e00000001,
104'h346b2191d60dbc631b00000000,
104'h2cf2be5ae5651711ca00000000,
104'h662da34f5b2432754800000000,
104'hb800308d0028ea195100000000,
104'h34be777a7c0eef5d1dffffffff,
104'h2878f6abf10c9bdf1900000000,
104'h08dff0bcbf48e2d79100000001,
104'h66b7963e6fe1397ac200000000,
104'h04bffa847ff80e5ef000000000,
104'h34ba8b94750c27cd18ffffffff,
104'hbc8b84fe1777012fee00000000,
104'h288895ba11b3ff6c6700000000,
104'h0486b1140dec1446d800000000,
104'hbc57c27dafa128b84200000000,
104'h2cd5bc72ab2a665f5400000000,
104'h00833a62066e37cddcf1722fe2,
104'h2ce2ad84c5d897f4b100000000,
104'h301bccbd37640885c800000000,
104'h660bbf79179947443200000000,
104'h2c9f3b963e1d9a7b3b00000000,
104'h54068e3b0db14c4a6200000000,
104'hb82247b944cfad0e9f00000000,
104'h602402734867b4c1cf00000000,
104'h28f97cb4f2d01b58a000000000,
104'h5460fd93c11b80273700000000,
104'h00acbcd059b8f8387165b508ca,
104'h94efc5c0dfcb1bb69600000000,
104'h08c18d1c83436a478600000001,
104'h28a631ec4c899e6a1300000000,
104'h08a8216250b647e06c00000001,
104'h907c95c1f91dc5013b6150c0c2,
104'h94d72830ae8473220800000000,
104'h00096dab12c6adf48dd01b9f9f,
104'h60e256d0c476f5e9ed00000000,
104'h04a5cad44be25582c400000000,
104'hb817b54f2f7eddcdfd00000000,
104'h34a67f2a4cf1d1a6e3ffffffff,
104'h60efaa78df0ad82f1500000000,
104'h30d6095aac374e1d6e00000000,
104'h2c5bc7d9b77c8e27f900000000,
104'h661b40cf36e9c860d300000000,
104'h66c055bc8019c0953300000000,
104'h66f8c1b2f1ba8bac7500000000,
104'hbc249f2f499524102a00000000,
104'h345118f5a2286cff5000000000,
104'h66e5fdfacb0afcf91500000000,
104'h309bb03e37dcc714b900000000,
104'h04f9a6aef30d7b691a00000000,
104'h667679ffec0e36671c00000000,
104'hbc893494121cd73d3900000000,
104'h30405d5f80a515324a00000000,
104'hbc75f5b9eba72c0e4e00000000,
104'h3428624b509db7743b00000000,
104'h600ef6e91d6c153fd800000000,
104'h28dd9d70bbe466e6c800000000,
104'h9405cfaf0be009e4c000000000,
104'h60cbdc3a97a71f084e00000000,
104'hbc6e2e59dceb78e0d600000000,
104'h009110d422d90912b26a19e6d4,
104'h005423efa821a4cb4375c8baeb,
104'hbc177e2d2e63b805c700000000,
104'h343530436a4b40019600000000,
104'h6080a3ec014224978400000000,
104'h00680ddbd0e0c89ec148d67a91,
104'h30ccea82998169460200000000,
104'h283f3e077ed0a47ea100000000,
104'h94ec0f18d8e33e50c600000000,
104'h347254d3e4acfd405900000000,
104'h2ca24f9a449e35b03c00000000,
104'h281a0509341d5c3f3a00000000,
104'h2c6e56b7dc77b723ef00000000,
104'h304aec35953006936000000000,
104'hbc5be7d7b733bc216700000000,
104'h541b1ea336e7191ace00000000,
104'h2c6f4b29de164beb2c00000000,
104'h289e73603c1d64753a00000000,
104'h601579952af2b778e500000000,
104'h2c2590394b9f08f83e00000000,
104'h54c508cc8a04958b0900000000,
104'h66cbb5b89711d2c52300000000,
104'hbcbbd736778e7e981c00000000,
104'h901f4b2b3e0955b312161e982c,
104'h9c8578020afa88e0f580080000,
104'h60712a9be262c963c500000000,
104'h00b65f1c6cf8845ef1aee37b5d,
104'hbc16acd72dc4a52e8900000000,
104'h3407cd2d0fd5f6ccab00000000,
104'h54aa756854ddfc30bb00000000,
104'h04c07ba2800bd7ab1700000000,
104'hbc17fe9f2fc199468300000000,
104'h941608ab2cbe0c307c00000000,
104'h34fde582fb78db0ff1ffffffff,
104'h30f3232ee6a8a35e5100000000,
104'h90b2f5e065aa4fe05418ba0031,
104'h044e76db9cb6d1ec6d00000000,
104'h60f9f646f3f011dae000000000,
104'h90fe581afc3fae597fc1f64383,
104'h9c3033ff6039e2d7733022d760,
104'h00b5301c6aa4acde4959dcfab3,
104'h6682cf1405570875ae00000000,
104'h9092a8cc25cddb7a9b5f73b6be,
104'h3076c657ed83e80e0700000000,
104'h947598d3ebbfdde87f00000000,
104'h08cfc34e9f9762be2e00000000,
104'h66faafa0f547a9a38f00000000,
104'h66a1a64a432bf1635700000000,
104'h54d3e15ca77801e9f000000000,
104'h2818d25331e08096c100000000,
104'h9ce492f6c974b3b3e96492b2c9,
104'h044539398a8d0cb81a00000000,
104'hb84e86199dc791be8f00000000,
104'h28f42782e806fddf0d00000000,
104'h085b8531b73b308b7600000000,
104'h9464d081c9d143eaa200000000,
104'h04efcf68dff7624eee00000000,
104'h28639a3fc7d43276a800000000,
104'h28f144ace25b7307b600000000,
104'h9018298730f91cdef2e13559c2,
104'h34cf51aa9ed22472a4ffffffff,
104'h90922de42445b23d8bd79fd9af,
104'h34179bcd2f9b6a0c3600000000,
104'h2ce0eda4c1d3196ea600000000,
104'hbcc36d3e8647e50f8f00000000,
104'h904191d583bccd1079fd5cc5fa,
104'h2ca9e0ee53622079c400000000,
104'h9cb0323e60e3377ec6a0323e40,
104'hb842ce8785818d020300000000,
104'h66e7a170cf1e0ed53c00000000,
104'h66a676744cc33d2a8600000000,
104'h949bf8b4373a70ef7400000000,
104'h9075ede3eb64612dc8118cce23,
104'h9c7be417f7e0bf68c160a400c1,
104'h08184abd30fa8304f500000000,
104'h0044ae65893e3b9d7c82ea0305,
104'h66788fb1f185826e0b00000000,
104'h28f50d28ea0e62ab1c00000000,
104'h66305829605750e5ae00000000,
104'h00eaacb0d560096bc04ab61c95,
104'h90cb4450968d6da61a4629f68c,
104'h00767c07ec32387b64a8b48350,
104'h9c8f25161e9821ac3088210410,
104'hb833b8f767c4c8368900000000,
104'h28f4e824e90b7bb51600000000,
104'h9c2dbc0f5b38bcbb7128bc0b51,
104'h2cbe43e87cb60c3a6c00000000,
104'h94a0849841dc61e2b800000000,
104'h6654238da8b9617a7200000000,
104'h66e004a0c03f274b7e00000000,
104'h00d9d2fcb320437140fa166df3,
104'h34b22cf464e93c4cd2ffffffff,
104'h3020eae7412eafd95d00000000,
104'h2c27b91f4f52ec09a500000000,
104'h0869fcb5d367962fcf00000000,
104'h00bfbb6c7f77b957ef3774c46e,
104'h349dfe943b0453ad08ffffffff,
104'h0461e8e9c3213ad54200000000,
104'h346c776fd859ef51b300000000,
104'h947ba55ff7c5b6de8b00000000,
104'h2c7a6af5f46815d9d000000000,
104'h284bcf5b97967f902c00000000,
104'h048e058c1c8dd5bc1b00000000,
104'hbc294c2b521a0ec73400000000,
104'h9c630867c6201b3b4020082340,
104'h045053dba06de21ddb00000000,
104'h0493f56c275dec4fbb00000000,
104'h90827d34040c16ed188e6bd91c,
104'hbcc3fb4c87fe64b2fc00000000,
104'h908589c40bb0c65661354f926a,
104'h66f5a170eb5471e7a800000000,
104'hb84cf1d799bb21327600000000,
104'h34ba340674c44f2488ffffffff,
104'h665a3079b4264c1f4c00000000,
104'h28a5eff84b06c1670d00000000,
104'h909fcf743ff5fb76eb6a3402d4,
104'h6034eef36976136bec00000000,
104'h54f33358e6b2cf566500000000,
104'h300cd3611960d1adc100000000,
104'h54d9276eb2526f9ba400000000,
104'h004734718e1e46693c657adaca,
104'h2c3929c572a767de4e00000000,
104'h9430ca0f6160b59bc100000000,
104'h084377238634c37d6900000000,
104'h9ca958e2520158ff020158e202,
104'h6695d7182b0169950200000000,
104'h9c105e5d20421c0f84001c0d00,
104'h946b27f3d6c738fe8e00000000,
104'h906a7ca9d441180b822b64a256,
104'h9461aabbc399e4583300000000,
104'h662ba6b15719cfeb3300000000,
104'h04240f3d48e18dfec300000000,
104'h66d20c20a4f02c6ee000000000,
104'h080140070245240d8a00000001,
104'h943dc5677be1380ec200000000,
104'h543eee637de07c5ec000000000,
104'h28713fabe2959b082b00000000,
104'h34b2de5c65e23090c4ffffffff,
104'hbc2668df4cf1d758e300000000,
104'h60eef2c2dd6d39fdda00000000,
104'h66649babc92044b94000000000,
104'h900bf91f175a4dc3b451b4dca3,
104'hbc034b7b06f0cca8e100000000,
104'hbcdf35bebe34f8bb6900000000,
104'h04c5707a8a4a66619400000000,
104'h0426afad4d907b822000000000,
104'hbc79b399f32a52e15400000000,
104'hbcf83cb4f09066762000000000,
104'h284b5a7f966d18e1da00000000,
104'h007f4d65fe40f5b381c043197f,
104'h342ff39b5f5d40dfba00000000,
104'h08d57906aa1b2d133600000001,
104'h041dc2173bc3d1168700000000,
104'h6081c9a603d0b432a100000000,
104'h9c76e9dfedf68984ed768984ed,
104'h60eac812d53b726d7600000000,
104'h34d55ba0aa1fdfe53fffffffff,
104'hbcc747d48e0ceae11900000000,
104'h662380c747bcbbb07900000000,
104'h6659f339b39958663200000000,
104'h60ada77c5b0bf2291700000000,
104'h6603974d07da899cb500000000,
104'hbc982eb030eb8244d700000000,
104'h00782fddf0867cde0cfeacbbfc,
104'h2ce6720ccc5f90c3bf00000000,
104'h90a2b37045d5bc48ab770f38ee,
104'hb8fe75fefcbf24207e00000000,
104'h9c039f59075579b7aa01191102,
104'h285553b1aa42a0978500000000,
104'hb81643a12ce16ac4c200000000,
104'h08b0650e60700421e000000001,
104'h5408cf1111a164cc4200000000,
104'h002730c74ea0e27e41c813458f,
104'hb8d31b3aa6a6b8ee4d00000000,
104'h90d21642a49e212a3c4c376898,
104'h28783865f08550020a00000000,
104'h66d1b9aea30d735f1a00000000,
104'hbcfeb99efd0486a70900000000,
104'h901b2ff9362c961b5937b9e26f,
104'h046bc0b3d7c3c9368700000000,
104'h9c34eacd69164c172c14480528,
104'h08ccca2e996eefcfdd00000001,
104'h66d06492a08d19d01a00000000,
104'h941c395d38de5a4abc00000000,
104'h94ec8c7ad907c1850f00000000,
104'h948ca448193ecc457d00000000,
104'h9cecf26ed97b7f2ff668722ed0,
104'h2c86dfc00d1d091d3a00000000,
104'h60d1b31ca320048b4000000000,
104'hbc66cb4fcdf12feae200000000,
104'h287c23eff82935135200000000,
104'hbcc2dd408585d78e0b00000000,
104'h60ac3f125832a2076500000000,
104'h08ca6ea09456eaa1ad00000001,
104'hbc22cf7145d8c65eb100000000,
104'h5406c73b0dc4437e8800000000,
104'h66145cbb28bc02d87800000000,
104'h288ae99c15b408446800000000,
104'hbcd8d756b1e959f0d200000000,
104'h945e1f11bc00c6cf0100000000,
104'hb88404740864ebe3c900000000,
104'hbcad43a25acf50b69e00000000,
104'h60d2aa00a55232aba400000000,
104'hb80ed2211da8575c5000000000,
104'h9c987aa230f5fe04eb907a0020,
104'h54e5b014cbf1c7d8e300000000,
104'h549ac1ca358e2f6c1c00000000,
104'h34aeb9ca5d23e70b47ffffffff,
104'h3083cfa407bb361c7600000000,
104'h94c50e508ad62d8aac00000000,
104'h345b251bb6f74b14ee00000000,
104'h90e91b72d27fe3b7ff96f8c52d,
104'h34ae5fd85c576d0daeffffffff,
104'h549669b82c887daa1000000000,
104'h2856e64bad921c822400000000,
104'h54f42872e803b7430700000000,
104'h0888539e1007d7b30f00000001,
104'hbcec79acd83570196a00000000,
104'h9c93a3c0274956999201028002,
104'hb8b67e2e6cb9478c7200000000,
104'h008b1f58165786efafe2a647c5,
104'h54df218abee9f8b6d300000000,
104'h28b307d8669948343200000000,
104'hbc9ca60639e47676c800000000,
104'h286b0367d642e7a58500000000,
104'h90f8f0b2f142c76585ba37d774,
104'h2cfc48f2f8ab5c385600000000,
104'h9c1e95593d6aa1dfd50a815915,
104'h28788c27f1cb42ae9600000000,
104'h60d4a286a90bc8011700000000,
104'h3095a9702be19982c300000000,
104'h30f52d86ea2a23a75400000000,
104'h943211fb64fa3cf0f400000000,
104'h046a9e65d5cfa26a9f00000000,
104'h94edf7b0dbd222f4a400000000,
104'h66ffbbeeff41d1ad8300000000,
104'h540539410a55574baa00000000,
104'h300e77af1c573a85ae00000000,
104'h60560e15acb2b76e6500000000,
104'h60d979f2b2487dd39000000000,
104'h5440725980c16e9a8200000000,
104'h9c1c6dc53819302f3218200530,
104'h54ca52fa943431cd6800000000,
104'h341f0cf13e7475f7e800000000,
104'h303479a568d63bc2ac00000000,
104'h0856ec05ad995f463200000000,
104'h34ec38c4d8ce08f49cffffffff,
104'h9c64064bc8b303fa6620024a40,
104'h6085d7840ba1d3a04300000000,
104'h9cf409cee8b85fac70b0098c60,
104'h2c2bbdd15779cfc3f300000000,
104'h94d8635eb0afedbc5f00000000,
104'h30ae60565cdc2714b800000000,
104'h665b0a85b6f30542e600000000,
104'h9c20ec8141deb516bd00a40001,
104'h669e0d8e3cccf51e9900000000,
104'h08aeb47a5d8a83001500000000,
104'h2c91dd842391dfe82300000000,
104'h66155b332aed03d2da00000000,
104'h30ce5a389c0957ff1200000000,
104'h54efc052df1310452600000000,
104'h345a9e31b5c8bb7c9100000000,
104'h08bdac487be9a2d4d300000001,
104'h082f8abd5fd9503cb200000000,
104'h54543c3fa8c053be8000000000,
104'h000113e902c61fde8cc733c78e,
104'h90230e2146e994fed3ca9adf95,
104'hb89a4c7e34ed93bcdb00000000,
104'h007a2c9df4b4ae50692edaee5d,
104'h28d8320ab0b2d0f06500000000,
104'hb8bcbb1c79bd792e7a00000000,
104'h2c0f38d91eead458d500000000,
104'h042c61cf584ddcd99b00000000,
104'h666797f7cfa14e924200000000,
104'h90b9799a724d0a479af473dde8,
104'h607c552ff8113ff72200000000,
104'h9403f83307f87838f000000000,
104'h0449110f926d54a3da00000000,
104'h60791bfdf2629f27c500000000,
104'h303292e165d40070a800000000,
104'h3039d8297373754fe600000000,
104'hb8b614b06c8b5b001600000000,
104'h603600a36ce6aaaccd00000000,
104'h280b4f4d1660bbadc100000000,
104'h00a836125083a4fa072bdb0c57,
104'h34c5463e8ac8158e90ffffffff,
104'h2cde91e8bd8b3bb81600000000,
104'hbc3dd3d57b1713852e00000000,
104'h30fc1250f817341f2e00000000,
104'h0457f519aff7f42cef00000000,
104'hbc1ec6353de77d2cce00000000,
104'h54e4d5d6c9f025dee000000000,
104'h3016b9412dd92b9ab200000000,
104'h54b79c9c6f96a2b82d00000000,
104'h30999fe0330335e70600000000,
104'h5433f6b567d60c94ac00000000,
104'h549f43423e34f04d6900000000,
104'h30e3642ac6568913ad00000000,
104'h0852ad53a55248c9a400000000,
104'h005d43cdbaeb5d8cd648a15a90,
104'h60c414b888c9c3169300000000,
104'h308d9f241ba04b1c4000000000,
104'h9c4788e78f2034b1400000a100,
104'h2c26b6814dc2aaa08500000000,
104'h662c5e03584e40d79c00000000,
104'h90c94ce8920248b504cb045d96,
104'h943958fd726b9481d700000000,
104'h302fb42f5f8601b60c00000000,
104'h30199b7f33e3e26cc700000000,
104'h546798d9cf901dbc2000000000,
104'h00a64ff64c319f1963d7ef0faf,
104'h30e68e36cd0e6ca91c00000000,
104'h00b9158e72da7cbcb493924b26,
104'h66055a550a3222156400000000,
104'h00f32c32e629a755531cd38839,
104'h042e01fd5ceb715cd600000000,
104'h54a560904ae3c0a0c700000000,
104'h30c894ba91e4e99ac900000000,
104'h60c4b81289f09c1ae100000000,
104'h34b2b8da655a91adb5ffffffff,
104'hbc97dce42fb6bafc6d00000000,
104'h04cdf76a9be8c42ed100000000,
104'h088949f412a488464900000001,
104'h30f0c834e12ecb7d5d00000000,
104'h084a36ed942354b14600000000,
104'h60465dc78ce13db2c200000000,
104'h5432443b64f012b8e000000000,
104'h94e9316ad2a818ac5000000000,
104'h6087e7080f95d29a2b00000000,
104'h94444f2d88e49e06c900000000,
104'h941d95433b85fe520b00000000,
104'h2c8761da0e3aef1b7500000000,
104'h9c6fb197df0a559d140a119514,
104'h04397eff727b6909f600000000,
104'h002f376f5e0ca9f3193be16277,
104'h90b6b2e66d47c0a98ff1724fe2,
104'h9ce526f6ca705a95e0600294c0,
104'h28244c9d488fde981f00000000,
104'h941ab11d3579907bf300000000,
104'h0427e9ed4fc27b348400000000,
104'hbc32238b647e3a63fc00000000,
104'h666d4365da4d7a999a00000000,
104'hbcdc94aeb9dcc8c8b900000000,
104'hbcc6b84e8dca08a09400000000,
104'h66d84fb2b0f4a9e8e900000000,
104'h66749ab7e9f074e8e000000000,
104'h04640083c89c85be3900000000,
104'h9cdf3b6abe2fcecb5f0f0a4a1e,
104'hbc929fcc25523a07a400000000,
104'hbccfb5f49f8541660a00000000,
104'hb86c1efbd820963d4100000000,
104'h28f37ca2e6ef2f94de00000000,
104'h2c86d43a0df6d79aed00000000,
104'h5436a47f6d980ff23000000000,
104'h5485a6740bede51edb00000000,
104'h6040f155819508dc2a00000000,
104'h08a6f95a4db74b866e00000001,
104'h3421a1b143d44c6ea800000000,
104'h9c505953a031f94b6310594320,
104'h00f5fae0eb9734842e8d2f6519,
104'h5442e78d85e0baa8c100000000,
104'h281694f12d941eba2800000000,
104'h2ce485f2c9be759c7c00000000,
104'h2c1766ab2e9c086a3800000000,
104'h60c9c33293ac25e05800000000,
104'h66a6919a4d5feab5bf00000000,
104'h306c86b7d97498f5e900000000,
104'h3415ee0d2bb1d6706300000000,
104'h66bb7cac7621ea134300000000,
104'h341b570f365dd03dbb00000000,
104'h08ee41fedc20be354100000001,
104'h0013b66b27766c75ec8a22e113,
104'hb8ca5058946d4019da00000000,
104'h34d4d0aea9b12b3462ffffffff,
104'h9044aa2789c5dc3a8b81761d02,
104'h00d9d124b32e94595d08657e10,
104'h042c4697589fbcd63f00000000,
104'h305695dbadca137c9400000000,
104'h34493d95925905e9b200000000,
104'h347dbb99fbcd93fa9b00000000,
104'h341cb3c939e4d12cc900000000,
104'h280569ef0aa4dcf24900000000,
104'h302d86a35becea1cd900000000,
104'hb8b6df286decad3cd900000000,
104'h908db84e1b2549f94aa8f1b751,
104'h0094bc5029f99776f38e53c71c,
104'hb8049bb7094d53b99a00000000,
104'h60e41132c8b29dfc6500000000,
104'hbc09c087131ad01d3500000000,
104'hb824285d485b8eebb700000000,
104'hb87c9f2df90aa99d1500000000,
104'hbcc1131882ab201c5600000000,
104'h94c504d08ad36876a600000000,
104'h340cf5731948cb2f9100000000,
104'h94c83f6490f56ea6ea00000000,
104'hb8cc1238988e697a1c00000000,
104'h9cdf0990bea4f3e64984018008,
104'h2c5f96f5bf2990215300000000,
104'h2cb836c07009c1b71300000000,
104'h085b27f5b6f8abf8f100000000,
104'h04d41f20a890af4e2100000000,
104'h2c112c43223fdda17f00000000,
104'h2804cb9f09caddae9500000000,
104'h0461d9abc31195752300000000,
104'h541ee1e53d16b38f2d00000000,
104'h90d900bab286ef900d5fef2abf,
104'h08c750608e0e996d1d00000001,
104'h94e698bccd23cfd14700000000,
104'h0809ba3d13797585f200000001,
104'h28be0bbc7c82bdd00500000000,
104'h2c23a3654738e7d37100000000,
104'h04284289502480eb4900000000,
104'h60b05c8660714613e200000000,
104'h085470aba8ff7c3efe00000000,
104'h6021af0d43e757bece00000000,
104'h9c73a06fe72acaa55522802545,
104'hbc314923624fd2179f00000000,
104'hbcaafee255c11aba8200000000,
104'h34b6e9b66d0c941319ffffffff,
104'h60a8e7d251d74adcae00000000,
104'h340f4c731e93a2702700000000,
104'h04e8b1c6d122c5274500000000,
104'h94ffd5c4ff7be3aff700000000,
104'h90713a0fe2ab9b7457daa17bb5,
104'h34c2fed685eb9c04d7ffffffff,
104'h669a30b634a663624c00000000,
104'h00a9819453e4a96ec98e2b031c,
104'h902424874851d24ba375f6cceb,
104'h907c44adf8aa7fac54d63b01ac,
104'h00af4f105e74194de823685e46,
104'h348b0788163de4397bffffffff,
104'h005d209bbad40140a83121dc62,
104'h2c13ce5527aa6a4c5400000000,
104'hbc288c3551c9c6c49300000000,
104'h606f0dffdea1aee84300000000,
104'h904113a982c3b6348782a59d05,
104'hbc2c983359a054c44000000000,
104'h34749385e95a87adb500000000,
104'h340d47591a98c05e3100000000,
104'hbc73cf13e7517b09a200000000,
104'h66856aa00adf93f2bf00000000,
104'h947dbc5ffb9e33e23c00000000,
104'h0033f1f567d5eb7cab09dd7212,
104'h08bd90367b54559ba800000001,
104'h2c7a5a03f48d58b81a00000000,
104'h34678a25cf10df492100000000,
104'h3021583542619f21c300000000,
104'h66608077c14147cd8200000000,
104'h34b646b86c442ff588ffffffff,
104'h60fc2c36f86259bfc400000000,
104'h940d50771a35662d6a00000000,
104'h281e35313c12cf7d2500000000,
104'h08145d21282782874f00000001,
104'h66c9fdf29395af222b00000000,
104'h94e2bd1cc547677f8e00000000,
104'h90ed2fc6da20668d40cd494b9a,
104'h90b1959a63671551ced680cbad,
104'h30f106b8e210a7552100000000,
104'hbc290c875205e5f90b00000000,
104'h305e5d97bce602dacc00000000,
104'h302e34895c3289336500000000,
104'h34a079ea409b463636ffffffff,
104'h941db9113b42c07b8500000000,
104'h54b2980065bb96487700000000,
104'h601f4a4b3e1cdb0b3900000000,
104'h084436e7884f4ba99e00000001,
104'h94fdc920fb8ef1e21d00000000,
104'h08a02468407c8eb5f900000001,
104'h28b0333e60efe3badf00000000,
104'h5462490fc477b389ef00000000,
104'h607f4f11fe0611110c00000000,
104'h04c83428901f56013e00000000,
104'hb87417c5e8efd820df00000000,
104'h9c2867c3506035b7c020258340,
104'h347ae947f589d0e61300000000,
104'h90dc64a4b83cd20b79e0b6afc1,
104'h04676c3fce8ec91c1d00000000,
104'h9ca976605214c6152900460000,
104'h54c5421e8a6d8043db00000000,
104'h08743f3de887e4b40f00000000,
104'h0021710d4290239220b1949f62,
104'h90cb04489611148322da10cbb4,
104'h94388ff971918a062300000000,
104'h6692b94e2534ebdd6900000000,
104'h0035b28d6b9c305c38d1e2e9a3,
104'h34e2ccdcc5e00cdec0ffffffff,
104'h00ee1536dceef510dddd0a47b9,
104'h04dbb43cb7514165a200000000,
104'h94c589208b43945f8700000000,
104'hb804377b08ab57085600000000,
104'h08a7a0364f92e4422500000000,
104'h04797d65f20abb2b1500000000,
104'h044199278372d079e500000000,
104'h30fdd784fbbad6e27500000000,
104'h04690b5bd20a167d1400000000,
104'h90b24e2864e72b10ce556538aa,
104'h605b52ffb655c189ab00000000,
104'hb806ec5b0de42c4cc800000000,
104'h2841bd01833c669b7800000000,
104'h002dcbe75bebdef4d719aadc32,
104'h3426730b4cab20705600000000,
104'h661ce15b39ea3324d400000000,
104'h9c46278b8cb84b827000038200,
104'h34ea8800d5b520b86affffffff,
104'hbc6a81abd588020e1000000000,
104'h0410cde521cc834a9900000000,
104'h94b94956726e5811dc00000000,
104'h30e37fd4c67db63bfb00000000,
104'h3424533d488b57421600000000,
104'h6644f55b8906f0a10d00000000,
104'h28662cc7ccdcbb24b900000000,
104'h28659cc5cb16615d2c00000000,
104'h283788216f816cee0200000000,
104'h2c1a471b34c10b068200000000,
104'h9c29683952aabfa05528282050,
104'h3415342f2acd5ffc9a00000000,
104'h34500cb9a0776bf3ee00000000,
104'h9c0dde871bed9e5adb0d9e021b,
104'h2caa9e0e55b44c626800000000,
104'h60a387724745ebfb8b00000000,
104'h34f39964e73ed92d7dffffffff,
104'h948682fe0d5a327db400000000,
104'h2c45fca78b85644c0a00000000,
104'h2c3443f5683fbb3b7f00000000,
104'h94c332828661157fc200000000,
104'h2c5227e1a4ae8b4e5d00000000,
104'h0825be634b45a63d8b00000001,
104'h2c73030fe64e7f979c00000000,
104'hb8eca874d982ddc60500000000,
104'h60d36c8ca65c28b1b800000000,
104'h548ba9a01713cd152700000000,
104'h3058ca25b18166f40200000000,
104'hbccc17989837cae76f00000000,
104'h60df1c64be7dc681fb00000000,
104'h944a90c395d12fb4a200000000,
104'h9ca18a9643fa9b2ef5a08a0641,
104'hb8bd684e7a45d1bd8b00000000,
104'h6049aec793a6dc9e4d00000000,
104'h906fd229df5d40fbba3292d265,
104'hbcf1a1c2e376c22bed00000000,
104'h001dcef93b58c329b1769222ec,
104'h3424c71549a31eec4600000000,
104'h901cd82f39410fc7825dd7e8bb,
104'h66ab590a56c47dc28800000000,
104'hb87d4bf7fa25cc0d4b00000000,
104'h60acb4ae5925fd4b4b00000000,
104'h5490993a21cac6fa9500000000,
104'h947465cde82bebdd5700000000,
104'h28002ba700fef548fd00000000,
104'h30e5f2f2cb6a2397d400000000,
104'h666117a7c2992d743200000000,
104'h046b696bd6c626528c00000000,
104'h00f08668e1d6a3baadc72a238e,
104'h90eaa940d5c0f9b0812a50f054,
104'h34e4e1d8c99726162effffffff,
104'h040d71431ac4c30a8900000000,
104'h087fc09fffb318446600000000,
104'h9ce82afad012237b2400227a00,
104'h60cc922c99672fbfce00000000,
104'h30cb76b696a953de5200000000,
104'h30b80aa87091efc42300000000,
104'h34cc777e984b00d396ffffffff,
104'h28ec4f02d83ee54f7d00000000,
104'h664fdf259f6ce6b5d900000000,
104'h549de0e43bbba31a7700000000,
104'h60a3ba2e47be2d9a7c00000000,
104'h08354abd6a327da76400000000,
104'h0073fbede79785662f0b815416,
104'h08818bb40387072a0e00000001,
104'hbca5ca6a4b7301b3e600000000,
104'h94df43b8bef04ba2e000000000,
104'h94e58a72cb47b5db8f00000000,
104'h9c809f76018cccce19808c4601,
104'h94f3ab90e76510f9ca00000000,
104'h30c2045884ec3e28d800000000,
104'h007c3411f829f9eb53a62dfd4b,
104'hb8377c8b6e4b00eb9600000000,
104'h28050d010ab3ab4c6700000000,
104'hbcdee2fabdfb6014f600000000,
104'h903f0e2b7e604f7bc05f4150be,
104'h54a2cf5245388c5f7100000000,
104'h9cc5ca1c8bc15c9082c1481082,
104'h281a4201345f5847be00000000,
104'h001a1a213459b06bb373ca8ce7,
104'h9031102f6248b4099179a426f3,
104'h66636a43c6436ca58600000000,
104'h60250fc94a41e9a18300000000,
104'h0043c5518799929833dd57e9ba,
104'h6004037d08de98cabd00000000,
104'h2ccaa0d495415f678200000000,
104'hb89646b42ca073004000000000,
104'h0052691da46f67e7dec1d10582,
104'h0862399dc430b7836100000000,
104'h00d4cd32a90474b708d941e9b1,
104'h04346d2368a76f484e00000000,
104'h0401cae3039e1e323c00000000,
104'h60588ef1b11c69113800000000,
104'h2c257abb4af72876ee00000000,
104'h2c6f1575de7df557fb00000000,
104'h00a89c0451f39f5ee79c3b6338,
104'h908babd817696257d2e2c98fc5,
104'hb8b7e0cc6f74b287e900000000,
104'h66085e091081380c0200000000,
104'h605df9e1bbd05148a000000000,
104'h2c3984b3737d3435fa00000000,
104'h301c62cb388886c41100000000,
104'hbcee7140dcf0064ae000000000,
104'h08ceedd89d9e95d23d00000000,
104'h906ad9e1d57ecb89fd14126828,
104'h2c661015cc9dd5103b00000000,
104'h9045057b8a064aed0c434f9686,
104'h30c3ed4a873a4adb7400000000,
104'h0854b7c1a9e9f134d300000000,
104'h04c82406901f094d3e00000000,
104'h549edd183d888cd81100000000,
104'h08565997ac484a439000000000,
104'h66e9f6b2d392ca162500000000,
104'h9ce38606c7054b590a01020002,
104'h60674679cebf6eea7e00000000,
104'h54d60020ac7de9e9fb00000000,
104'h609cbb183919570f3200000000,
104'hbcc449708857ff13af00000000,
104'h2c7b9bfdf7e33002c600000000,
104'h085e9a43bdd87baeb000000000,
104'h304ff5539fccf5009900000000,
104'h308f2da41e9c445a3800000000,
104'h30f4c404e9f72b02ee00000000,
104'h661d4d613ac4cd728900000000,
104'h3478e1bff1ffdcc6ff00000000,
104'h08df1e04be3477136800000001,
104'hbc20b0ed411556c92a00000000,
104'h04462adb8c36a9176d00000000,
104'h007088bde1caa344953b2c0276,
104'h08d2b1f0a5afaf1a5f00000000,
104'hb8abe11a5729c6375300000000,
104'h9cb9b00e73b0547860b0100860,
104'h00f53eaeea3fb95b7f34f80a69,
104'h60c9acc4930940511200000000,
104'h04fadee8f51e282b3c00000000,
104'h9c5a465fb43a117b741a005b34,
104'h94dc23f4b80eebe71d00000000,
104'h34d27de6a4d83a94b0ffffffff,
104'h28b3c0bc67754787ea00000000,
104'h3411c32923499dfb9300000000,
104'h2cf2a4ece598e3ca3100000000,
104'h94c7c0b28f6ee9c9dd00000000,
104'h2877a8f3ef568b2bad00000000,
104'h0486e7ce0d99b3da3300000000,
104'h300ff9f71f72a5e5e500000000,
104'h661dbc893bea55ccd400000000,
104'h90cc45ea980975f512c5301f8a,
104'h2c82e1ae05f188f8e300000000,
104'h3456a777ad591315b200000000,
104'h905fe4cbbf31c27f636e26b4dc,
104'h603552076ae126c4c200000000,
104'h6606ca2b0ddc4f36b800000000,
104'hb8a5fdc64b94683c2800000000,
104'h045e58d9bce62fbecc00000000,
104'h287e13a5fc97d87c2f00000000,
104'h601126a12250b473a100000000,
104'h9c3b994b77cbbe3c970b980817,
104'h940b64111641d96f8300000000,
104'hbc32dd27651a61fb3400000000,
104'h081368732648628f9000000001,
104'h9c84e262094889f39100806201,
104'h6008fdd311e7b76ecf00000000,
104'h2c4a8ceb95c3b6208700000000,
104'h04176cff2e477f698e00000000,
104'h60208d6d41aa1c405400000000,
104'h60e64980cca2fd9c4500000000,
104'h34000d53000863cd1000000000,
104'h3094fda429d42ce2a800000000,
104'hb8101ac9200922051200000000,
104'h080d16791a169bd92d00000001,
104'h90dbd4bcb79215e02449c15c93,
104'h60f74fc8eede08dabc00000000,
104'h9c1956d9328b241e1609041812,
104'h305f601dbe5cbe05b900000000,
104'h08ed658adacb133c9600000000,
104'h90d284c4a515ad332bc729f78e,
104'h9057d9fdaf660773cc31de8e63,
104'h6084cdcc09964c002c00000000,
104'h0434ce1b69d9bebcb300000000,
104'hbcc929fc92342fc96800000000,
104'h54fe8892fd538cdba700000000,
104'hbce832e6d06a69abd400000000,
104'h903c28cf780c174718303f8860,
104'h3021b8d14332a27f6500000000,
104'h664912fb9274d13be900000000,
104'h66650ecbca75f6e3eb00000000,
104'h08e11c04c2b337b66600000000,
104'h000c169f18719333e37da9d2fb,
104'h089d75983aa5cd724b00000001,
104'h34a50cda4aab0f8a56ffffffff,
104'h544e5a1f9c6ed6eddd00000000,
104'h049714c82ed08bc6a100000000,
104'hbcdd78c6ba40d6618100000000,
104'hbc2d84755ba08b804100000000,
104'h3425217b4ae8c7cad100000000,
104'h9455f0adabb592186b00000000,
104'h04e830e8d0521ce7a400000000,
104'h541cf8fb39d17ea6a200000000,
104'h34d6bc7aad00792f00ffffffff,
104'hbcb5d3ac6b04a80b0900000000,
104'h544b7e5f963b2de37600000000,
104'h009899cc31ccb8dc996552a8ca,
104'h2c2e017d5c6675fbcc00000000,
104'h0403532706074b7b0e00000000,
104'h28258d874bc672348c00000000,
104'h30e9c248d3544601a800000000,
104'h9008d2e311a7e50c4faf37ef5e,
104'hbc1ff07d3f43f64b8700000000,
104'h083656c16caaaebe5500000000,
104'hbc4b79cf966cedf3d900000000,
104'h30419f0d83aa09465400000000,
104'h04e7990ccf459e598b00000000,
104'h04211e6f427e8461fd00000000,
104'hb867f3c1cf5db495bb00000000,
104'h54c8e0569195c1882b00000000,
104'h544626378c533587a600000000,
104'h60ddf4f0bb1beff93700000000,
104'hb8860f7c0c9f59c63e00000000,
104'h94ee9d26dd3308b16600000000,
104'h28fcdd5ef91729b32e00000000,
104'h085b36a5b673ca69e700000001,
104'h2c66d865cdbbd9667700000000,
104'h08dbe7d6b7b4759e6800000000,
104'h2817efdf2f36e4bf6d00000000,
104'h544f0beb9ed1488ea200000000,
104'h30d305d8a61deb553b00000000,
104'h663c5ecd78f2bb34e500000000,
104'h3413fb1b27da4c88b400000000,
104'hb838e925718d7b4a1a00000000,
104'h90d87b36b0d08372a108f84411,
104'h0417ac652f1828513000000000,
104'h90b38872672342f34690ca8121,
104'h60930eb22632cf816500000000,
104'h60b7c7de6f2e51a15c00000000,
104'h34db06feb6bc27d478ffffffff,
104'h28848d44099525da2a00000000,
104'hbc3408f368108e0b2100000000,
104'h3481a732038141bc02ffffffff,
104'h2c92b0fc256ec09fdd00000000,
104'h3415eaf32b6c4f23d800000000,
104'h28e03046c03e5bcd7c00000000,
104'h2c648091c991fba62300000000,
104'h905378bda6b4159068e76d2dce,
104'h28dceedab9e594a8cb00000000,
104'h000b290d160fb9a71f1ae2b435,
104'h60a9e75a532763414e00000000,
104'h00d438a0a86fe58bdf441e2c87,
104'h60cad25e9575c84feb00000000,
104'h08c963a492f78476ef00000001,
104'hbc641af1c876186bec00000000,
104'h2c3757076ec10b688200000000,
104'h66923adc24f137f2e200000000,
104'h2cf19c70e3db751eb600000000,
104'h00cb86b0977ff703ff4b7db496,
104'h00044651084cfe1199514462a1,
104'h909cb9b639a32d76463f94c07f,
104'h006e5bd1dcd7a07caf45fc4e8b,
104'h004c41fb986396e9c7afd8e55f,
104'h285104dda2fb505ef600000000,
104'h94b04c4a60556eb9aa00000000,
104'h66bf76227e71f771e300000000,
104'h30439031879bcbfe3700000000,
104'h281b9d0d372131334200000000,
104'h9044dbfb8947bd9b8f03666006,
104'h28ab8bc6573dc6dd7b00000000,
104'h906d60b1da2f26255e42469484,
104'h34d3a53ea71ceb6f39ffffffff,
104'h3489be24131757fb2effffffff,
104'h6021891f43ef37a0de00000000,
104'h0001cedd03cf71389ed14015a1,
104'h6013bfd5276165f1c200000000,
104'hb81b3429369677b82c00000000,
104'h084a268b94dece9abd00000000,
104'h0482a21405e9351ad200000000,
104'h308b1b2c16f1a39ae300000000,
104'h6667eb6bcf93d2b82700000000,
104'h2cc9686892fcecacf900000000,
104'h9c38cdb771a335ac462005a440,
104'h3416f1a92d4c434b9800000000,
104'hb8c67d448c921ad42400000000,
104'hbc301f1b60354eb56a00000000,
104'h6061f123c3cdf2ce9b00000000,
104'h540c09a718c6ffe28d00000000,
104'h603aef1b756f7df3de00000000,
104'h289d66fe3a428d958500000000,
104'h660dd7bb1bc3285e8600000000,
104'h30b03588605a3043b400000000,
104'h54ec324cd8fd25ecfa00000000,
104'h9c90287420f19e2ae390082020,
104'h94abf8dc57354e3d6a00000000,
104'h2ce3d3aec7dc4748b800000000,
104'h0049a4399386b8a80dd05ce1a0,
104'h04e897ded1d55156aa00000000,
104'h9c48f7eb91ef184ade48104a90,
104'h60fb4e74f6ad53d45a00000000,
104'h28e08e40c149d8019300000000,
104'h9419b59d3369d3fbd300000000,
104'hb87c2445f882f6680500000000,
104'hbcc89c4091d280c8a500000000,
104'h04e1a5c2c3dda1dabb00000000,
104'h908ace0c15a82ef65022e0fa45,
104'hbc04f94909ea9474d500000000,
104'h60d4bf6ca98195020300000000,
104'h08568c21ad8a30101400000000,
104'h9c28f98f5109c7291308c10911,
104'h90189e5731165a4f2c0ec4181d,
104'h00c9465e921c736538e5b9c3ca,
104'h30074eb90e9018882000000000,
104'h90289c8551fbdd72f7d341f7a6,
104'h085f66d1be6cebd9d900000001,
104'h6009cb73139c9acc3900000000,
104'hb80fe6ed1f5fed1dbf00000000,
104'hbcf6e74eedc30eb28600000000,
104'hb8a25214443aa8f17500000000,
104'h907d7509fa6ea61ddd13d31427,
104'h9c25ba1b4bc1bbb28301ba1203,
104'h345b564bb6ced3c89d00000000,
104'h04288b8551112d792200000000,
104'h9c88758210bdcc347b88440010,
104'h308d19a21aec8e24d900000000,
104'h28c931da927d0199fa00000000,
104'h54c4ea808916d1512d00000000,
104'h28358b3f6b2f5ff15e00000000,
104'h66bec2e87d8dea581b00000000,
104'h90e10e5cc24d48fd9aac46a158,
104'h28937266264628578c00000000,
104'hbc8f809e1f0e50371c00000000,
104'hb8bd5f467ac152288200000000,
104'h00224c314484b6d809a703094d,
104'h9066d297cd9d826a3bfb50fdf6,
104'h302aac0155e6a7e2cd00000000,
104'hb81b042136f7c378ef00000000,
104'hbccc97b89941340d8200000000,
104'h28e5e672cb3e6b6f7c00000000,
104'h00de6fc6bc910dd4226f7d9ade,
104'h00aeb2d65dcf38289e7deafefb,
104'hbcf16954e2fd0576fa00000000,
104'h08593559b27d2b43fa00000001,
104'h60aeba4e5dae44ee5c00000000,
104'h34f9d8c6f3da2616b4ffffffff,
104'hbcb585626b824bf80400000000,
104'hbc2872ab50e045c4c000000000,
104'h66e585facb92ac0e2500000000,
104'hbc3dcf537b56ff25ad00000000,
104'h60c27c42844e84719d00000000,
104'h9c07fdc90f0ffad51f07f8c10f,
104'h545c5929b8a1be164300000000,
104'h90415bd982d7b130af96eae92d,
104'hb8e82a56d06607bfcc00000000,
104'h28d66210acb5c6546b00000000,
104'h54f5c63aeb1991e53300000000,
104'h28c62fba8cd9261cb200000000,
104'h66ee37fedc978ac42f00000000,
104'h9429d6e3534be0259700000000,
104'hb846eb8f8d4e5a5b9c00000000,
104'h08ae68565c4ac3c79500000001,
104'h2c9599982b2f9e635f00000000,
104'h308dbfa01bdcbc22b900000000,
104'h9c70f387e155e659ab50e201a1,
104'h00d20f0ea405ec110bd7fb1faf,
104'h34ca0f86941c2f7738ffffffff,
104'h30702babe0b28a2e6500000000,
104'hbc2a9481552320bb4600000000,
104'hbc84994009357cd96a00000000,
104'h0803a627078006e20000000000,
104'h94bf565c7ef6b62aed00000000,
104'hbcf990def31190672300000000,
104'h30ca684c94ad50005a00000000,
104'h60d835d8b0b649846c00000000,
104'h6037271d6e4167f78200000000,
104'h549c36fe38e0d838c100000000,
104'h003e49977c31bb67637004fedf,
104'h08bce2fe79c5f83c8b00000001,
104'h665eb147bd1903713200000000,
104'h04a2e142452037114000000000,
104'h54a6f6784daf10ec5e00000000,
104'hb8f79df8ef456fef8a00000000,
104'h0435b43b6b61a879c300000000,
104'h3439760b720a07d11400000000,
104'h303c945779611e71c200000000,
104'h9cc0a32481ade9745b80a12401,
104'h66921b5a24bcb2f07900000000,
104'h0820e7b341cf41569e00000000,
104'h049e34903ceaadd4d500000000,
104'h9093fae2271ef9b33d8d03511a,
104'h342d7e075ad83ab8b000000000,
104'h66d8b4a0b152f685a500000000,
104'h94775485ee5d04f7ba00000000,
104'h28b2f994659211882400000000,
104'h60629f9bc5ae93ae5d00000000,
104'h2cf8672ef055d639ab00000000,
104'h28d55d94aa2f65b95e00000000,
104'h00d5bf9aab7dfdd5fb53bd70a6,
104'h289aef7c35b5cdb26b00000000,
104'h54b915c27211ab552300000000,
104'h542d251f5a268df94d00000000,
104'hbc0cb95319ea6778d400000000,
104'h046c0909d8ff34a6fe00000000,
104'h28aee2b85d44dcb98900000000,
104'hb8106c85202c37995800000000,
104'h90d21f1ca4f35352e6214c4e42,
104'h6065339fca46d06b8d00000000,
104'hb8b27c7064aded425b00000000,
104'h9c936124261698772d12002424,
104'h904b755d96bca24279f7d71fef,
104'h088ce2a019f2e4dce500000001,
104'h00fa9d4cf5f6fbd2edf1991fe2,
104'h28621c61c45fe275bf00000000,
104'h08bb0c6c76d5912aab00000001,
104'h2c8e356e1c0371dd0600000000,
104'h34658babcb11434b2200000000,
104'hbc8623960ccdc3709b00000000,
104'h662180b1430c38eb1800000000,
104'h669677662cf1b34ce300000000,
104'h34f299ece5009a8901ffffffff,
104'h04dbe828b708e54d1100000000,
104'h900f3a891eb10e6062be34e97c,
104'hb8e29fe8c57fa10dff00000000,
104'h606ba671d716f46f2d00000000,
104'h3438477570246de74800000000,
104'hb8a5ee524b4a626f9400000000,
104'h66fcd256f9776efbee00000000,
104'hbc3e9b997d9fdfda3f00000000,
104'h2c3e0adb7c157f212a00000000,
104'h60ca1c6e94b7e1f26f00000000,
104'h2ca9de0e535b0cf7b600000000,
104'h2886efc20dfc07aef800000000,
104'h04e367bec61ab6d93500000000,
104'h2884913e09c615cc8c00000000,
104'h9486be720d03a6e30700000000,
104'h044725518e2cb2cb5900000000,
104'h90a77f7a4e13aef127b4d18b69,
104'h9093e5222731e2e163a207c344,
104'h94561ae3ac31249f6200000000,
104'hb8d24aa0a4cf440a9e00000000,
104'h9077df73efc87d4690bfa2357f,
104'h902dfc795b1c0a093831f67063,
104'h04fdc6bcfb09aa091300000000,
104'h94657a15ca88ba541100000000,
104'h904601078c2133bd426732bace,
104'h2cf187a0e3eca828d900000000,
104'hbc344161688917001200000000,
104'h94f15a0ae2e13084c200000000,
104'hb84cc995994d60319a00000000,
104'h540782ff0fa6b6204d00000000,
104'hbcde3630bce08768c100000000,
104'h60139ce5278f5d7a1e00000000,
104'h60060a7f0cdb8c84b700000000,
104'h9474b6ede9ab88ce5700000000,
104'h541bfc8b37c5d31e8b00000000,
104'h00408101813414196874951ae9,
104'h30d00122a0c0be968100000000,
104'h009b37ce36ee5114dc8988e312,
104'h660717d10eb30e046600000000,
104'h901c50c13885c33c0b9993fd33,
104'h0042d6e3854ff8499f92cf2d24,
104'hbcebe604d7979bd02f00000000,
104'h901fb7633f1607fb2c09b09813,
104'h0004e28309ebf5c8d7f0d84be0,
104'h9436211d6c21b7794300000000,
104'h66c7edec8f18d1e33100000000,
104'h086a369fd46fccdfdf00000001,
104'h90cb18a8968ad29a1541ca3283,
104'h30766133eceb7608d600000000,
104'h289247e624afb82c5f00000000,
104'h303c9ce579642491c800000000,
104'h009c619238be9c947d5afe26b5,
104'hbc2a8483554729d78e00000000,
104'h90f13854e259ef8fb3a8d7db51,
104'h00bc1d9678b912f272753088ea,
104'h081c379d380732970e00000000,
104'h90e9646cd26ac4c5d583a0a907,
104'h043fcf977f3874e77000000000,
104'h300a9813154657e58c00000000,
104'h04ada12c5b638f7fc700000000,
104'h947f4655fecfb4b09f00000000,
104'h602f6a0b5e632117c600000000,
104'h902417bb48d4ef44a9f0f8ffe1,
104'h94ecb09cd91d4a2d3a00000000,
104'hbc635b95c6ca637c9400000000,
104'h2c993010322c28fd5800000000,
104'h306c53efd8ee90f2dd00000000,
104'h00580453b0041583085c19d6b8,
104'h60dd4190ba11b7072300000000,
104'h947f960bffd39d78a700000000,
104'h9cec300cd89d30d03a8c300018,
104'h942a46ab5419405f3200000000,
104'h9cda81a8b53691316d12812025,
104'h903fdc597faaeb6e559537372a,
104'h603f3b757e1a7ebf3400000000,
104'h6063ae05c7ab35a25600000000,
104'h3074113be80b4fd91600000000,
104'h94f38f58e7a85bb85000000000,
104'h04313189626f669bde00000000,
104'h9c037cc306e0fc2cc1007c0000,
104'h2c23d1a947fb4ce0f600000000,
104'hb802076d046a933bd500000000,
104'h600b79a7160390450700000000,
104'h60718143e3b5b6de6b00000000,
104'h08aa105054525e27a400000001,
104'h94e1e8f2c3ac12d45800000000,
104'h9c92a730251cdf9f3910871021,
104'h901795e72f642499c873b17ee7,
104'h08a306944674558de800000001,
104'h9c0aa44b1526b7654d02a44105,
104'h60b3f986674ef4899d00000000,
104'h602b210d564220378400000000,
104'hbccc59d2980480f10900000000,
104'h2815f5d72be739ccce00000000,
104'h9ce2dc06c5daaae0b5c2880085,
104'h04a695164d0c209f1800000000,
104'h54fa9b6cf5fd2a34fa00000000,
104'h341165f72210aeeb2100000000,
104'h602666114cfd9a86fb00000000,
104'h0872f063e5a0b8ac4100000000,
104'h9cbec8c07db717366eb600006c,
104'h00ffc908ff10079f200fd0a81f,
104'h00d6db06ad31975d6308726410,
104'h28c13d52822c17415800000000,
104'hb8bbcb3077e109d8c200000000,
104'hb88abf6c153f90cb7f00000000,
104'h940b2a47165c3143b800000000,
104'h2c94124428c3873c8700000000,
104'h04abf81a57673ff9ce00000000,
104'h9ce43584c8fa734ef4e03104c0,
104'h94b66f326cee3416dc00000000,
104'h5479119bf270ef7fe100000000,
104'h301690df2d4af3779500000000,
104'h08d7e3b0af2034094000000001,
104'h3075712beaf327b8e600000000,
104'h347269b3e4ae52e85c00000000,
104'h60b542e06a69da37d300000000,
104'hb80cce4f190833db1000000000,
104'h340c238d1810d00b2100000000,
104'h9c1054ef20515059a210504920,
104'h2889a77a1335a6136b00000000,
104'h0876c5c1ede52fa2ca00000000,
104'hb89325b82676aceded00000000,
104'h60ba99ac75e6a2b0cd00000000,
104'h90a2c410455b84f1b7f940e1f2,
104'h30f7e664ef98c0423100000000,
104'h28554311aabd7a3c7a00000000,
104'h082a0a4f547da0d1fb00000001,
104'h60928a02255ba0abb700000000,
104'h6032189b64f6da98ed00000000,
104'h085cf2f3b9b6afda6d00000000,
104'hbc12053524e3bd96c700000000,
104'h949356ae26109f272100000000,
104'hb88890c411794f85f200000000,
104'hbcb1d8c0632c01a95800000000,
104'hbcf9f4baf35007e3a000000000,
104'h345d7377ba27223f4e00000000,
104'h08514f43a2634be9c600000001,
104'h284643db8c8edf861d00000000,
104'h2c46cf478d7eaa97fd00000000,
104'h28ac95b8598547d80a00000000,
104'h3036a0736d54d8a5a900000000,
104'h5494af9e2997f5522f00000000,
104'h30749733e93c6c917800000000,
104'hbc755ed7eaa229ce4400000000,
104'hb8c89cb4914e5a979c00000000,
104'h2ced436cdad6aaecad00000000,
104'h287fdae5ff6230b3c400000000,
104'h34cadc2e95cd5e069affffffff,
104'h603ea86b7d2412a14800000000,
104'h307352a7e630a4376100000000,
104'h547f34b9fe4075db8000000000,
104'h2c740723e866765bcc00000000,
104'h9c68f3f5d1619da1c36091a1c1,
104'h60cadcaa9551410fa200000000,
104'h906ccb0fd97ad6ebf5161de42c,
104'h04314511620480b10900000000,
104'h00d1fbb0a39d74763a6f7026dd,
104'h60760cdbec091d571200000000,
104'h301fd0493f538ac3a700000000,
104'hbcb1e758638d86e21b00000000,
104'h60100801203c6c077800000000,
104'h2ce2ba96c59d90ee3b00000000,
104'h547602c5ec66e43fcd00000000,
104'hbc39ab5f733e0ed77c00000000,
104'hb846ad438da5352a4a00000000,
104'h2827e93d4f082fb51000000000,
104'h54ad2ce45ad6d244ad00000000,
104'h60f63a7ceca09a664100000000,
104'hbcd84bd6b0e3dcc6c700000000,
104'h2873482de62649894c00000000,
104'h28eca506d9e65fb0cc00000000,
104'h3004aa1709752777ea00000000,
104'h2847901f8fbd4bba7a00000000,
104'h6626b2c94dd86a4cb000000000,
104'h2cfecd8cfd0533630a00000000,
104'hbc26fb8d4d88afe61100000000,
104'h2848f27b9132c6e56500000000,
104'h66a5b06e4b11d9e12300000000,
104'hb83a94d5754b103d9600000000,
104'h94299c3d537ca995f900000000,
104'h2c04374908756f27ea00000000,
104'h90d2f480a5d81c22b00ae8a215,
104'h549cf5403963551dc600000000,
104'h28f8e588f17e8663fd00000000,
104'h0085eee80b49c15f93cfb0479e,
104'h003dde5f7b3270f364704f52df,
104'h5412752f24e87ce4d000000000,
104'h90669ccfcdef342ede89a8e113,
104'h3460f5bdc1db166cb600000000,
104'hb8fff966ff0954331200000000,
104'h08f0a700e12f9e735f00000001,
104'h669f73703efa9cdaf500000000,
104'h547ff425ffff2332fe00000000,
104'h044a7cf994f5fdc2eb00000000,
104'h089fa9143f83eca80700000000,
104'h545086cda11f26453e00000000,
104'hb826de7f4de97890d200000000,
104'h28a3cc764701e1810300000000,
104'h0073a5cde7d23666a445dc348b,
104'h087ce045f9a5324e4a00000000,
104'h9424752d484f03659e00000000,
104'h94d4f740a9562f4dac00000000,
104'h28b653866cc466888800000000,
104'h9c02f53705069ed70d02941705,
104'h3033c48d67f98c90f300000000,
104'h548738b20edb5308b600000000,
104'h08e074a4c04d03f59a00000001,
104'hbcd22702a44645bf8c00000000,
104'h308da4fe1bcb38f29600000000,
104'h3091783222c874949000000000,
104'h2c03578506a2b1864500000000,
104'h9cd0430ca0377ce56e10400420,
104'h08aa3ae45432096b6400000001,
104'h66f5c91ceb22f7cf4500000000,
104'h34625689c4abae1e5700000000,
104'h046f02afdeb5962a6b00000000,
104'h9432769f640b5add1600000000,
104'h348eead01d2dfc975bffffffff,
104'h003c581178d9549eb215acb02a,
104'h94f18b4ce3cb5f6e9600000000,
104'h9c21948b43f76622ee21040242,
104'h946dc8b1dbc9dece9300000000,
104'h54c54e788a739be5e700000000,
104'hbc61ee47c3caa2929500000000,
104'h60169d092d1cc0213900000000,
104'h2ce6fa1ccdc3b6568700000000,
104'h604fb8279f5496d3a900000000,
104'h2836a8fb6d53a575a700000000,
104'h90d5e47aab5bd9b7b78e3dcd1c,
104'h94504271a014d70d2900000000,
104'h54a61f744c13f4472700000000,
104'h08a824ca504ca9f79900000001,
104'h66fa8b40f5f27fc2e400000000,
104'hbc6e1113dc1250d12400000000,
104'h90949ac829a27f224436e5ea6d,
104'h28b637146cc96df69200000000,
104'h54d7fdb8af8f5b261e00000000,
104'h9491015e228c6f841800000000,
104'h04a24c7e44559e47ab00000000,
104'h66dda13abbe2ab56c500000000,
104'h348b744216d570c0aaffffffff,
104'h30635ab5c6de3b08bc00000000,
104'h34fae2f6f562d491c5ffffffff,
104'hb87d909bfb7d97f5fb00000000,
104'h603d73437a4fa1719f00000000,
104'hbc669077cdecf73ad900000000,
104'h3488189210cb40e096ffffffff,
104'hbced1e96da0365b30600000000,
104'hbc934b1226d42a18a800000000,
104'hb820c2054117a3fb2f00000000,
104'h343b33b176b71e186e00000000,
104'h3040d08d8108c26f1100000000,
104'h90509817a1582399b008bb8e11,
104'h28fa3abcf4167d2b2c00000000,
104'h308686b20d4143178200000000,
104'h08c017de80e5580aca00000001,
104'h9c28c2af513302cf6620028f40,
104'h28caf1fe95ca7aaa9400000000,
104'hb806eff70db2a2bc6500000000,
104'h540ad1eb153b4c657600000000,
104'h90c07f3880d2189ca41267a424,
104'h60180b2d30fcd058f900000000,
104'h045d59dfba2dcbe95b00000000,
104'h66eec810dd6ec15fdd00000000,
104'h30df4e14bedc11e0b800000000,
104'h340155a5020e6e151c00000000,
104'h04383ac970ca697c9400000000,
104'h94ed2fb4da0d54d71a00000000,
104'h54d0fba4a1c4777a8800000000,
104'h9cdeccc8bd977fc02e964cc02c,
104'h308d15161a20c2594100000000,
104'h90702a31e025a0af4b558a9eab,
104'h30f72048eecf2e4e9e00000000,
104'h008e17f81cf6ed3ced85053509,
104'h9c01f727034539598a01310102,
104'h60b044e8608ebac41d00000000,
104'h2c8aa05e1583f7360700000000,
104'h04700a93e0d1da66a300000000,
104'h2886fb5a0d33cd636700000000,
104'h0849f93d931fb4fb3f00000000,
104'hbc8d2c461a91ef162300000000,
104'h281623f72c83271e0600000000,
104'hb81fc8113fab99525700000000,
104'h60832c8a06d71d2eae00000000,
104'h2ceac064d5230ecf4600000000,
104'h60a00f86407aef47f500000000,
104'h90dd0faaba7a5409f4a75ba34e,
104'h3040b03581f27d42e400000000,
104'h08cb2512969fab3c3f00000000,
104'h28c924a0928e0abc1c00000000,
104'h040610870c37d0676f00000000,
104'h54abc19857f5db14eb00000000,
104'h28136eb526e1f542c300000000,
104'hb8a5e6a64b358d636b00000000,
104'h2c721507e4717d4be200000000,
104'h28878a180fa338864600000000,
104'h28177dab2ed979beb200000000,
104'hb81184f923be47187c00000000,
104'h9c11f3892345e5978b01e18103,
104'h90369f136de21376c4d48c65a9,
104'h047b7e53f69ea1903d00000000,
104'h08cb5af4966843bdd000000001,
104'h54a98e6e53703029e000000000,
104'h347081e9e196e5c62d00000000,
104'h6645690d8af6319aec00000000,
104'h60446ffb88764b2fec00000000,
104'h30b9541872c39fe28700000000,
104'h94a71ff84e6aa555d500000000,
104'h2c1e823b3d44cabd8900000000,
104'h901cf76d392d61515a31963c63,
104'h9097bee22f1713a52e80ad4701,
104'h041c52a3388244020400000000,
104'hb8c4da3c89f269d4e400000000,
104'h2851d0a9a3c446028800000000,
104'h9cbad53275a0864c41a0840041,
104'h60a75f4a4e262faf4c00000000,
104'h04accd70593de7c57b00000000,
104'h661a07113442f5238500000000,
104'h0031a96363c08eba81f2381de4,
104'h602a774b5459d23bb300000000,
104'h54d28436a580796a0000000000,
104'h9c745205e8522691a4500201a0,
104'h604dd9d99b3ddfd17b00000000,
104'h66b8380670631185c600000000,
104'h90bb72f076e12fa6c25a5d56b4,
104'h346494e3c9face2ef500000000,
104'h307d10f1faf0c86ce100000000,
104'h30692adfd241cf6f8300000000,
104'h90a7d9fe4f78775df0dfaea3bf,
104'hbce15f0ac2559bddab00000000,
104'h6652850ba5deb370bd00000000,
104'h9ce14530c21769d72e01411002,
104'h54f445bee8e39966c700000000,
104'hb8716bdfe22a7b795400000000,
104'h34c0788880c5a7ba8bffffffff,
104'h3485685e0a7e3a9ffcffffffff,
104'hbcab0e9256483aa99000000000,
104'h287922bdf28014e20000000000,
104'h0481b9c80317c82d2f00000000,
104'hb860e1c7c1d117a4a200000000,
104'h0845d8d98bc7dc028f00000000,
104'h30381707701b4bfd3600000000,
104'h04b3232c6666d3a7cd00000000,
104'h08baeaca7562d2cbc500000001,
104'h9c9f14f03e635a53c603105006,
104'h2876881dedeec0a6dd00000000,
104'h089d1b123a3fa5057f00000001,
104'h305c28c9b8a5b9ee4b00000000,
104'h9c137f3d264e6e7b9c026e3904,
104'h00e2e15cc57a4ebff45d301cb9,
104'hb8ad13dc5a75b32deb00000000,
104'h30842d22084316f38600000000,
104'h04d3a01ca7b32d586600000000,
104'h281f3a273e1a8e253500000000,
104'h609f0be83ede90fabd00000000,
104'h908ef5361d22afb545ac5a8358,
104'hb8654befcae587cccb00000000,
104'h2c7ed5ddfd4852bb9000000000,
104'h28d70d98ae7d6d4ffa00000000,
104'h2c4a6a6794624617c400000000,
104'h66552313aa06cab90d00000000,
104'h0073a3dde7c82c60903bd03e77,
104'h30eaaf4ad51e930b3d00000000,
104'h60fbe210f73d17f77a00000000,
104'h281811eb30191efd3200000000,
104'h90abbf8857c9e6f49362597cc4,
104'h085a9361b562e90dc500000001,
104'h54159d952be35f34c600000000,
104'h041cd0d7398309760600000000,
104'h30def040bdf80a56f000000000,
104'h287be839f73b72377600000000,
104'h549c4a563841d1b58300000000,
104'h9c0d64351a02eb090500600100,
104'h284c296398775a69ee00000000,
104'h9c91e83423d4cd66a990c82421,
104'h543c81b179b921507200000000,
104'h54409c67811280912500000000,
104'h60e70a4eced6570aac00000000,
104'h081759b32ef2b57ee500000000,
104'h3410490720c57bee8a00000000,
104'h605b95cbb7ba62f07400000000,
104'h00355e676aecbc1ad9221a8243,
104'hbc380f1570bb815e7700000000,
104'h281491b929960b682c00000000,
104'h002338c146d58706abf8bfc7f1,
104'h34dc9d08b9ab017856ffffffff,
104'h347a66bbf4f3a3e4e700000000,
104'h344eb9259d9475a42800000000,
104'h347db9abfbc4bdb28900000000,
104'h08df6996bed9db06b300000000,
104'h0098cb0031a92bf05241f6f083,
104'h54a208ac44dc5c7cb800000000,
104'h04a418e8489233d62400000000,
104'h9c8b137016c9b8a49389102012,
104'h908b324c164f44659ec4762988,
104'h005535afaaa2ddd645f81385ef,
104'hbc83a2d80784f2520900000000,
104'h301515f52af24630e400000000,
104'h94c09ef88149b41f9300000000,
104'hbc47e18d8f8e138c1c00000000,
104'h004f6fdb9e245e054873cde0e6,
104'hbce89882d181eb8a0300000000,
104'h00889f6a11e85e00d070fd6ae1,
104'h30d819a4b0fc9384f900000000,
104'h9041e45183abb7ce57ea539fd4,
104'hbca3ee7c47dd4c94ba00000000,
104'h60accdfe59d2c0e8a500000000,
104'h9077d759ef3cef99794b38c096,
104'h9c8e309a1ced9c8edb8c108a18,
104'h90c617408c0ec92d1dc8de6d91,
104'h663a511574e377b8c600000000,
104'h9cf28006e5b535ae6ab0000660,
104'h9c81d11603a785244f81810403,
104'h040c3e311825fd354b00000000,
104'h907b5b0ff673b951e708e25e11,
104'h0062650fc4fa6fa0f45cd4b0b8,
104'h08d60e26ac4546758a00000001,
104'h087f3aadfe87408c0e00000000,
104'h9420aa4b4116d88d2d00000000,
104'h04d643d4acd82354b000000000,
104'h2c317c29621491592900000000,
104'h08311013622b27135600000000,
104'h669b092a36c5c4528b00000000,
104'h00a6c5b24d47d2a58fee9857dc,
104'hb8d97b7cb2e872b4d000000000,
104'h66aa6dc254ce00a69c00000000,
104'h60a4ce0c497a877ff500000000,
104'h907c000df8587b75b0247b7848,
104'h3493b884272cd36959ffffffff,
104'h34082f1f100f592b1e00000000,
104'h2cfb5b52f63bc8f17700000000,
104'h5402f443050617a50c00000000,
104'h30b7aba06f69f853d300000000,
104'h08c8db849181787e0200000000,
104'h34489f5b91984b8a3000000000,
104'hbc530fb3a6011d130200000000,
104'h0870192fe03802557000000000,
104'h904a265794a8e28051e2c4d7c5,
104'h003c948779926e2a24cf02b19d,
104'h9003abbf0765fda1cb66561ecc,
104'h282c918f59a26e4c4400000000,
104'h00f66ef4ecebd710d7e24605c3,
104'h34d6c134adfbabb2f7ffffffff,
104'h04f18dc4e364a72dc900000000,
104'h6642f12385fb951af700000000,
104'h9c2240bd4471d211e320401140,
104'h34dfb7c6bf401b0180ffffffff,
104'h2cb4672668d80398b000000000,
104'h66c0e04a81202ba14000000000,
104'h0099d30e33f30b60e68cde6f19,
104'h5492969a25a1eef64300000000,
104'h28c4554288cd78c29a00000000,
104'h606d5365da2ac2bf5500000000,
104'h00de894cbd77f6dfef56802cac,
104'h60768813ede4f674c900000000,
104'h944f617b9efc688cf800000000,
104'hbcfa0ad2f49747522e00000000,
104'h941472d72808c46b1100000000,
104'hb868428dd06a1c57d400000000,
104'h2cbf012c7e2db0d55b00000000,
104'h306512f3cad6823ead00000000,
104'h089fcb083f4cdfe79900000001,
104'hbcd3886aa7bae7827500000000,
104'h9ced95b8db932b7c2681013802,
104'h088a442414519861a300000001,
104'h34727949e41a71333400000000,
104'hb81ca80b3984fad40900000000,
104'h300bec83170f2e631e00000000,
104'h66e4c2cac9dd8a98bb00000000,
104'h040990f313f5dc2ceb00000000,
104'hb839fbcf7305952d0b00000000,
104'h6636bee56d6c0b69d800000000,
104'h54807f44009eb5ca3d00000000,
104'h301ad167358140b40200000000,
104'h047d6a17fae5116cca00000000,
104'h66bc32427883906c0700000000,
104'h041bb5f1375c52d1b800000000,
104'h54f22606e4dbfaacb700000000,
104'h2c8de53e1b8266720400000000,
104'h541157fd22568751ad00000000,
104'h34786f2ff043f68f8700000000,
104'h347f2633fef221f4e400000000,
104'h3090ebac21aea7205d00000000,
104'h3077ad71ef1435f32800000000,
104'h04ddff60bb1d11e53a00000000,
104'h6612954725bc0a6a7800000000,
104'h948407ba08d88254b100000000,
104'h30529c01a511de352300000000,
104'h28ca86e695ec71b0d800000000,
104'h30cbe2a8976dc3efdb00000000,
104'h04c64fce8ca7c2f04f00000000,
104'h542cf90b59b23df46400000000,
104'h90d4721ea807bed50fd3cccba7,
104'h30b6a9b46d969a622d00000000,
104'hbcd1e644a308cfd51100000000,
104'h306e85f1dd3d0f157a00000000,
104'h00bbf9687798fe2e3154f796a8,
104'h089831ca303095a76100000001,
104'h0025797d4aa82bde50cda55b9a,
104'h2cc1701082a687724d00000000,
104'h34aca1285992109e24ffffffff,
104'hbc6cee4dd99ff9983f00000000,
104'h9c5dc3d9bbddf5eebb5dc1c8bb,
104'h0427d0cd4f46d8f18d00000000,
104'h30aeb9b85d1033072000000000,
104'h9495fe9a2ba2c6184500000000,
104'h667f0bb7fe0968e71200000000,
104'hb8c12d828281b16c0300000000,
104'hbc48df7d912f7e475e00000000,
104'h9cb6ae126d3037096030260060,
104'h946ea379dd5c5ba5b800000000,
104'h663ff7957f5dbac9bb00000000,
104'hbc517ad5a24e673d9c00000000,
104'h0041f41583484449908a385f13,
104'h2c9c697c3816c10b2d00000000,
104'h940f0c611e0c1ae31800000000,
104'h04f0401ee0c13eca8200000000,
104'h04b7f4026fb321b66600000000,
104'h30dc4824b83227f76400000000,
104'h282735474e5ff39dbf00000000,
104'h00cfafba9ff5b1ceebc561898a,
104'h04937d3a26b0bf326100000000,
104'h2c6fb5cfdf7d3b4bfa00000000,
104'h9c94a7aa2935e2d56b14a28029,
104'h2c7e960bfd0649290c00000000,
104'h28e78b1ecf98489e3000000000,
104'hb83f34dd7e2741e74e00000000,
104'h30ac84e659cb826c9700000000,
104'h2c018b6f03bde9bc7b00000000,
104'h28acc50e5967a5dbcf00000000,
104'h9443d3ad87bb9ea67700000000,
104'h30f25a5ee406e8430d00000000,
104'h54947444280b54651600000000,
104'hb8befe687d42fac58500000000,
104'h2820aca1418d50701a00000000,
104'h54ada1725bae26385c00000000,
104'hbc9c00ec38e4a604c900000000,
104'h088ab68c15e4273cc800000001,
104'h04ec6616d89272202400000000,
104'h082f3f815e8eca2c1d00000000,
104'h34c72dca8e9ad77c35ffffffff,
104'h286a98ddd5fa4724f400000000,
104'h542ab27155afba965f00000000,
104'hb8c705ea8e955e002a00000000,
104'h3060c339c19d3daa3a00000000,
104'hbcb4fcb66979325bf200000000,
104'h66f5d00ceb73fcb5e700000000,
104'h5469320fd2d4e792a900000000,
104'h30d0d59aa1ad09705a00000000,
104'h9079657df2d8fcc0b1a199bd43,
104'h2858094db043a7598700000000,
104'h2803ed4f077e68c5fc00000000,
104'h304e45519c80c7ac0100000000,
104'h66ee028edc4576378a00000000,
104'hbcd5348eaaf44564e800000000,
104'h0484cd0809c85f749000000000,
104'h08c03eb880d7e13eaf00000001,
104'h348d2f4a1abdaa9a7bffffffff,
104'h5424343548d7fdb6af00000000,
104'h948e529e1cc645848c00000000,
104'h28cfba329ffe1b08fc00000000,
104'hbce2f310c52361cd4600000000,
104'h9418769f303913317200000000,
104'h54dd6b6eba3010d36000000000,
104'h6628fc2151bf15ea7e00000000,
104'h040a8143153a9faf7500000000,
104'h00bb7628764564b38a00dadc00,
104'h005ef0d9bd19b3413378a41af0,
104'h9ced14e2dac9cec293c904c292,
104'h00dbb93eb79924203274dd5ee9,
104'h309639382c69ed1bd300000000,
104'hbcf52840ea9a9aac3500000000,
104'hb85360d7a6841e720800000000,
104'h94c8a6669185eb000b00000000,
104'h9c2ad229551e43493c0a420914,
104'h34ed4300da6530f9caffffffff,
104'h9c7b085df64e39d99c4a085994,
104'h946b001bd6c8ac2e9100000000,
104'h349ddf5e3b201a1f40ffffffff,
104'h0424de7d494e5c039c00000000,
104'h086c7fd7d83631d56c00000000,
104'h66c1a9b883695b8dd200000000,
104'h34900b36201ec07b3dffffffff,
104'h00df8414bfc4fdac89a481c148,
104'h544b07a5961b734b3600000000,
104'h601e32a13c5fa8fbbf00000000,
104'h08278c114fd6a13ead00000000,
104'h944c2927983973d57200000000,
104'hbcb62c246c4247158400000000,
104'hbcc25634843280576500000000,
104'h3049a44f939cc3483900000000,
104'hb8baaf147575185dea00000000,
104'h9c5b45b9b6575217ae534011a6,
104'h082d7bd35a8789800f00000000,
104'h0404224f085a497bb400000000,
104'h9081633c02e1c122c360a21ec1,
104'h28b6f8be6de31530c600000000,
104'h901a36dd34a2a85a45b89e8771,
104'h2c26e0734df7f2b4ef00000000,
104'h00927f0024c140088253bf08a6,
104'h6006b5970d2d6d415a00000000,
104'h662bc6b357d57cc4aa00000000,
104'hb80d45191a3999d37300000000,
104'h94c1a7be8354e2eda900000000,
104'h046a38a3d49113282200000000,
104'h284b96b397dee29cbd00000000,
104'h6097c2a22f09b5bb1300000000,
104'h2cb96ed872f4f3b0e900000000,
104'h9c350a436a3f1bc77e350a436a,
104'h28b6be3c6d3a71c37400000000,
104'h6655576faa34d9496900000000,
104'h00a0d1ac4118383330b909df71,
104'h546ffed5df7277fbe400000000,
104'h00bb80b2775ffe19bf1b7ecc36,
104'h2cdd0ddeba95335c2a00000000,
104'hbc70b99de14b72559600000000,
104'h2c8ab6b8151374a72600000000,
104'h2c26cd734df3177ee600000000,
104'h00577c51aeae0ed85c058b2a0a,
104'h2cf97c06f218dff53100000000,
104'h943d1e517acb3aaa9600000000,
104'h2c61bfdfc3e289d2c500000000,
104'h2c38452770b7529a6e00000000,
104'h28985a4a30dfbaf2bf00000000,
104'h9098edfc31874ee40e1fa3183f,
104'h003f1f577e77dcf5efb6fc4d6d,
104'h042796bf4f1901853200000000,
104'h2c9d01cc3a9bb9323700000000,
104'h304b2a1b966d1237da00000000,
104'h3078df39f156d4c7ad00000000,
104'h541bab7b3756ba75ad00000000,
104'h9c5f0be7be9c8c8e391c088638,
104'h940da30d1b3d417f7a00000000,
104'h28dd9ee4bb6cf129d900000000,
104'h04a249b8446b384dd600000000,
104'h08037dfd062d62ed5a00000001,
104'h304875319027759f4e00000000,
104'h9c2e29bd5cd0edf8a10029b800,
104'hb85a43dbb493d1ec2700000000,
104'h2cf2496ee42c66275800000000,
104'h9ce388e6c70da3751b01806403,
104'h9caaf71e559243162482431604,
104'h049cf840398bfa321700000000,
104'h94fbcb9af7923c222400000000,
104'h6648129190379be16f00000000,
104'h9451aa6da378a465f100000000,
104'h9457d147af38bfff7100000000,
104'h082e4de35ce986bad300000000,
104'h0492128e24768bc5ed00000000,
104'hbcca930695b381c26700000000,
104'h3015c5532bc44e328800000000,
104'h2c5b85a5b7b663d46c00000000,
104'h00f1d53ee3b87c0070aa513f53,
104'h2c062c4b0c79870ff300000000,
104'hbc38d6bf71296bad5200000000,
104'h2c4e14439ccded4a9b00000000,
104'h303d73017a0bd1731700000000,
104'h2c8a9d9815981c283000000000,
104'h606393f1c72efb4f5d00000000,
104'hbcaf071a5e9db9023b00000000,
104'h66b250366412ccfd2500000000,
104'h00713a53e2f2e4f2e5641f46c7,
104'hb812974525d37bf6a600000000,
104'h049b578e366358d7c600000000,
104'h30e69d40cde70b7cce00000000,
104'h281401d728f3414ae600000000,
104'hbc66071bcc2888875100000000,
104'h04e96afcd253daada700000000,
104'h00ead67cd56d05d3da57dc50af,
104'h2c6b1f87d6e7cd12cf00000000,
104'h341b15d5369e57de3c00000000,
104'h281e92c53db3485e6600000000,
104'h049b444c361790e32f00000000,
104'h081a6ac33453e02ba700000001,
104'h2cb581d06bbf3cda7e00000000,
104'h66148c4b29dc27d2b800000000,
104'h00217b0f421b5d87363cd89678,
104'h042ee6e95d2f0e715e00000000,
104'h30d91570b25b2661b600000000,
104'h344f00e99e36fae36d00000000,
104'h04a5db224b1278a32400000000,
104'h288c43581814a7c52900000000,
104'h2cd32712a6231f4d4600000000,
104'h9c0106030221bf734301060302,
104'h603110eb620fcb171f00000000,
104'h9c0a5b7514633809c602180104,
104'h08541919a8b4ce7e6900000000,
104'h04c29cf885c76f628e00000000,
104'h34bd94c67b2299c145ffffffff,
104'h2842b69b854c071d9800000000,
104'h0858d9e1b115f6d92b00000000,
104'h2cf63328ece78090cf00000000,
104'h28792b15f24a05839400000000,
104'h340e082d1cd298dea500000000,
104'h9c4463cd889ff7383f04630808,
104'h2cde21f4bc8d64de1a00000000,
104'h943664356cd88b3ab100000000,
104'h54b1af8a63bc2d2e7800000000,
104'h60293d3b525b4a81b600000000,
104'h34622ebbc4b80a2a7000000000,
104'h280e1c891c4783c98f00000000,
104'h66bd38127a6f3fefde00000000,
104'h6642f88d85cb078e9600000000,
104'h94850adc0af15a56e200000000,
104'h9c30fc71617aa40ff530a40161,
104'h3097d9242fc308fe8600000000,
104'h949fb4203f2861455000000000,
104'hbc89d3b813d5bb40ab00000000,
104'h9ce8f84ad1737cede6607848c0,
104'h08bdf6227bbefc3c7d00000001,
104'h9cf99a58f30e26831c08020010,
104'hbcc992b0938b8eca1700000000,
104'h30cad0789574fb41e900000000,
104'h90ae9e6c5d4a498994e4d7e5c9,
104'h28c06192809442242800000000,
104'h9c38bd23712ab2d35528b00351,
104'h2c1791592f96e7ec2d00000000,
104'h90890d5e12cb5cc49642519a84,
104'h9452cc31a5db3b10b600000000,
104'h669cb46e3914013b2800000000,
104'hbc4e134b9cc967ce9200000000,
104'h085a2a5fb4b75dd06e00000000,
104'hbc682891d007b4230f00000000,
104'h007145f9e238cfe171aa15db53,
104'h00ec7ab0d8487bc79034f67868,
104'h281a08c93411b08b2300000000,
104'h30a9d11453adec3a5b00000000,
104'hbc7e2b1bfc5270a7a400000000,
104'h6061b7ebc37f80b9ff00000000,
104'h2c5967fdb2db74d2b600000000,
104'h907cac1df9ad3e3a5ad19227a3,
104'hb81c89393909b16b1300000000,
104'h902f07575e5caf7fb973a828e7,
104'h089f335c3e73068be600000001,
104'h2cfaac04f57ba101f700000000,
104'h902c71b3580e5c0f1c222dbc44,
104'h9c39715572149cfd2910105520,
104'h90760249ece37d92c6957fdb2a,
104'h281c4f3338e1276ec200000000,
104'h30ba61e6741eb6713d00000000,
104'h904b4a479655ba13ab1ef0543d,
104'h3429981d53242dc94800000000,
104'hb8122001242380634700000000,
104'h9c54c337a9ff0272fe540232a8,
104'h28c5b28c8bebd39ed700000000,
104'h2c34643f6848270d9000000000,
104'h00ce34d49ca176be426fab92de,
104'h9c116b012260fdf3c100690100,
104'hb882168404d39282a700000000,
104'h005d020bba9db5403bfab74bf5,
104'h28bdb00a7bde7162bc00000000,
104'h90431aa786bb62d276f87875f0,
104'hb8e3ae8ec7bdfb9c7b00000000,
104'h0483b8e007bde0447b00000000,
104'hbcb2400264fdf32cfb00000000,
104'h08deff86bd1166f12200000001,
104'h6018ff0f3103efcd0700000000,
104'h941ffc233f8bebf61700000000,
104'h60fb9f1ef7af1afc5e00000000,
104'h2892330224aa3c2e5400000000,
104'h668d585e1a09abf51300000000,
104'h046deb31db24d8374900000000,
104'h60b113bc628823b41000000000,
104'h00873a780eb8906a713fcae27f,
104'h2c8a56e2141248f52400000000,
104'h284bd16997bee0e67d00000000,
104'h942af03f55d1e432a300000000,
104'h04db874ab7f20d86e400000000,
104'h540962fb12833baa0600000000,
104'h9cc7a62a8f78fde7f140a42281,
104'h9cac130258c34f588680030000,
104'h54c4f6d68916d9612d00000000,
104'h60b531046a97d4f82f00000000,
104'h285c8cd9b91a63153400000000,
104'h663b666b762cf4055900000000,
104'h5467527dce6915dbd200000000,
104'h541b41613684c1bc0900000000,
104'hb8e054d0c0c200508400000000,
104'h04ad60d45a947d182800000000,
104'h5459cfa1b31460d32800000000,
104'h340d60711a0b8ad71700000000,
104'h3420f9754186017c0c00000000,
104'h54dd84a2bbc031748000000000,
104'h60dc8f9cb985542a0a00000000,
104'h54332695667e152bfc00000000,
104'h5432222564034e790600000000,
104'h6617e0332fb273f46400000000,
104'h28be1fd47cb105c06200000000,
104'h54cb782a963221936400000000,
104'h666aa23fd5dd0b22ba00000000,
104'h08b28de66515437f2a00000001,
104'h9cf0f9a8e14c87779940812081,
104'h669e05923c64ccf3c900000000,
104'h5411f923232c175b5800000000,
104'h00d7341cae15baef2becef0bd9,
104'h04d10276a2f4672ae800000000,
104'h941ccb31398e102a1c00000000,
104'h04bdd2327bde8f02bd00000000,
104'h087c8537f9af91245f00000000,
104'h04190ba132442ebf8800000000,
104'h54b5915e6b2440194800000000,
104'h9c5f84cdbf0749f90e0700c90e,
104'hbc8fbf921f689903d100000000,
104'h6088528410dde410bb00000000,
104'h54536c81a6cf8d9e9f00000000,
104'h00019453031d5c1f3a1ef0723d,
104'h084e2d939c7c4167f800000001,
104'h6038008570618903c300000000,
104'h28103cf7200d859b1b00000000,
104'h003530256a2b95555760c57ac1,
104'h60cea5949d771533ee00000000,
104'h30a0aafe41549b73a900000000,
104'h04162f1f2c4490ed8900000000,
104'h542fb3a15ff00178e000000000,
104'h90bb09fa76423b4584f932bff2,
104'h604fd3559ff99542f300000000,
104'h60b13b58624774778e00000000,
104'h5498262630eb686ad600000000,
104'h2c39c925739ef67e3d00000000,
104'h944d66e59a176c512e00000000,
104'h5490a6062148d1199100000000,
104'h6604bb190960ce0dc100000000,
104'h34075d6f0e1225c12400000000,
104'h54313f0f62b1127e6200000000,
104'h34387f89703ea3b17d00000000,
104'h942851d55044f23f8900000000,
104'h30bfcd3e7f3fc3e97f00000000,
104'h30e8a136d1acf5aa5900000000,
104'h94a3243c46b5c5206b00000000,
104'h00aff5bc5f1dd0df3bcdc69b9a,
104'hb8582aefb0b667d66c00000000,
104'h2c2bbeb7576c7fb7d800000000,
104'h2812bc8325156a472a00000000,
104'h00d05e30a0d221cca4a27ffd44,
104'h28c814e4902ac46d5500000000,
104'h04a334f246539681a700000000,
104'h0412bcbd2552a403a500000000,
104'h94836e8e0668d8ebd100000000,
104'h30e3357cc62328894600000000,
104'h66bd8d4a7b401beb8000000000,
104'h60a9654a5213df392700000000,
104'h0875b637ebb8a6187100000000,
104'h6662c317c512ff0d2500000000,
104'h0434bd1d69f16dd2e200000000,
104'h30b9428a724464c38800000000,
104'h04a3f08a470775350e00000000,
104'h041f00153ee64ed6cc00000000,
104'hb843a5cb875fe61bbf00000000,
104'h9092acde2517d9852f85755b0a,
104'h54a884e85199ee1e3300000000,
104'h2c78bad5f1fd3ac8fa00000000,
104'hb88b94b217045aa10800000000,
104'hbcb548a46a7dbe5ffb00000000,
104'h60b906b27232f4b96500000000,
104'h04f2cdb8e59781c22f00000000,
104'h66a9c336530f9d471f00000000,
104'hbcc1863c8304f02f0900000000,
104'h0053b549a78328e206d6de2bad,
104'h54fb9f1ef7affea05f00000000,
104'h947cd6b5f991fbea2300000000,
104'h289a2208342f27d75e00000000,
104'h909cfc083988667a10149a7229,
104'h9ce6a168cd4828499040204880,
104'h081a608f3492c06e2500000000,
104'h30b5a4686b347a356800000000,
104'h9c6cf253d9dd4560ba4c404098,
104'h6615d2f52b2391974700000000,
104'h60745e23e817b0b12f00000000,
104'h349fe1ba3f36d8296dffffffff,
104'h900cdb8919f89976f1f442ffe8,
104'h34533e25a6f3696ae600000000,
104'h08aeb8d25d1c8e933900000001,
104'h2cab7a5e56e58e94cb00000000,
104'h04a4a708495cf29db900000000,
104'h005a7957b4f1faa6e34c73fe97,
104'h3024c5fd497a97f3f500000000,
104'h60d35ab6a690c6582100000000,
104'h28587035b0b81cb07000000000,
104'h609226ec24ee2c28dc00000000,
104'h281ec7013dc006b08000000000,
104'h2ccc3b2298ad04525a00000000,
104'h3415fe6d2bf29f92e500000000,
104'h9cf57544eac700d28ec500408a,
104'hb83769436ef790b0ef00000000,
104'h604620018cc6a9648d00000000,
104'h3012450f242f3f255e00000000,
104'h042d9ec15b571783ae00000000,
104'h9c71461de25fe7cdbf51460da2,
104'h945dd9b3bbe5726cca00000000,
104'h04f6e37aedba7b467400000000,
104'h2cdb69beb6d02b1aa000000000,
104'h34fc62f2f81339eb26ffffffff,
104'h083e84977d5ff84dbf00000001,
104'h9cbfa5127fea0fd6d4aa051254,
104'h9c10a8a12186927a0d00802001,
104'h90abb124579eb0e43d3501c06a,
104'h00f3090ce61f2fe33e1238f024,
104'h6048013590ec74b4d800000000,
104'h30f9b9c6f32cc0815900000000,
104'h541a8e113589f2a01300000000,
104'h28679b77cf51ea0fa300000000,
104'h28889b4211885dc21000000000,
104'h28b7078c6e7ec40dfd00000000,
104'h9c82431804cea0f89d82001804,
104'h289b3c34369053b22000000000,
104'h3084c29c09cc3ae09800000000,
104'h54668859cd5dc801bb00000000,
104'h943f859b7f3fd9d37f00000000,
104'h340137a5026f75afde00000000,
104'h30e7f2a0cfadb7ec5b00000000,
104'h2c5d3e85ba5b933bb700000000,
104'h0007f6f90fe1b708c3e9ae01d2,
104'h3012a6272584b4e00900000000,
104'h305352afa6993cc63200000000,
104'h9490b87621b6089c6c00000000,
104'h66cfa4909f30ce816100000000,
104'h280fec1d1fd9522ab200000000,
104'h665b3629b6f16d50e200000000,
104'h6630908b61c2a7048500000000,
104'h005e87c5bd59b215b3b839db70,
104'h2cf239e6e4cdea6a9b00000000,
104'hbc349c6d697ea969fd00000000,
104'h606fed21dfca09549400000000,
104'h669605f22c606fabc000000000,
104'h608d0be21a6df681db00000000,
104'h2c12b0dd25ce8cf09d00000000,
104'h2c7f009bfe53666da600000000,
104'h0066707bcc38111d709e81993c,
104'h34dfaa72bf334b5166ffffffff,
104'h94344ad968836fc80600000000,
104'h34b4895669e01128c0ffffffff,
104'h007484c1e9ca1c50943ea1127d,
104'h5496a9f42d3999b57300000000,
104'hb8a16dbe4293e5ce2700000000,
104'hb8e751b6ce16f86f2d00000000,
104'h9c6eec1fddee1320dc6e0000dc,
104'h00bd6ac87ae1ee90c39f59593d,
104'h6098c8ee317a3ee3f400000000,
104'h08f7b018ef60271bc000000001,
104'hbc13bbf92750f371a100000000,
104'h309f99503fe632c4cc00000000,
104'h08ad37ca5a5406e7a800000001,
104'h668906de12f0440ce000000000,
104'h60e5f5aecb4cb7219900000000,
104'h04daadecb5dcab2eb900000000,
104'h349341b026f185bae3ffffffff,
104'h30eb4466d64412278800000000,
104'h6693069e26afd40e5f00000000,
104'h909f6cfa3e2b78b156b4144b68,
104'h309e9a023dd53f3caa00000000,
104'h2c346313680bf0471700000000,
104'h2808482b1074bc1de900000000,
104'h082366db466c1829d800000001,
104'h94efa020df23734d4600000000,
104'h3089e9401387594e0e00000000,
104'h66387fb170695d29d200000000,
104'hbc4277ef843ee2777d00000000,
104'hbc50df69a1819dcc0300000000,
104'h9c9a69523450641da010601020,
104'h08915e9222c6a1148d00000001,
104'h9c504897a08e8c7c1d00081400,
104'h00c48f3a89e5f69ccbaa85d754,
104'hb84701a78e9743922e00000000,
104'h5421022f42b7edbe6f00000000,
104'h9c19cd313343a71b8701851103,
104'h08c212f88456f19bad00000001,
104'h947cdc9ff9cdc6909b00000000,
104'h286b73e7d6d2a508a500000000,
104'h3016c61f2d681f2fd000000000,
104'h54237a03469abea63500000000,
104'hb83eb0997dc2d7f28500000000,
104'h66f02918e07da4d1fb00000000,
104'h08cb3fbe96babd9a7500000000,
104'h54c2ffb485d6c9a2ad00000000,
104'h60de3ff6bc2dfe9f5b00000000,
104'h545f8325bf48c6f99100000000,
104'h2c591271b2b2a73c6500000000,
104'h60c88b74911f3a6f3e00000000,
104'hb865d917cbaadd705500000000,
104'hbc804f6e0034615f6800000000,
104'hbc41629782f2dcf4e500000000,
104'h08a7309e4ef674e8ec00000001,
104'h2831d65b6324b3494900000000,
104'h34c547508ae8c5e4d1ffffffff,
104'h2c562091ac2dbba75b00000000,
104'h08caae9295bc98f07900000000,
104'h04ba1e2274b1db086300000000,
104'h3092902e25ddc268bb00000000,
104'h94db88bcb7787c2df000000000,
104'h08f4f0b2e90f02691e00000001,
104'h668ba2ca17df4b8ebe00000000,
104'h34333b69667220cde400000000,
104'h9cd9a37ab30eb36b1d08a36a11,
104'h344b8e5f9717c9312f00000000,
104'h9471e2b9e36c17bdd800000000,
104'h947ec65dfdf326eee600000000,
104'h349dc52c3b85d2400bffffffff,
104'h94154af32acd41269a00000000,
104'h00d06846a074ee71e94556b889,
104'h942e9a6d5d9416b02800000000,
104'h606c0e33d870a58de100000000,
104'h042795d54f217a2b4200000000,
104'h342c49db580f9a8d1f00000000,
104'h9ce38cf6c755adf1ab418cf083,
104'hb860eaebc172d631e500000000,
104'h94040a610821c01f4300000000,
104'h08e5a9d0cb5682f1ad00000001,
104'h54db5f5cb6dda690bb00000000,
104'hb88293b405c4690a8800000000,
104'h54a5eff64b061ae30c00000000,
104'h2c21368942e42a7ac800000000,
104'h94563efdac3e366f7c00000000,
104'h9c028cf505253efb4a000cf100,
104'h08ffb9f8ff30ce556100000001,
104'h60e1aa64c3beb00a7d00000000,
104'h90ac453858ad8f6c5b01ca5403,
104'h34af27045e4094e381ffffffff,
104'h542887c7511dda553b00000000,
104'h04514bc3a2b34e826600000000,
104'h6612f76f252d5f695a00000000,
104'h6094fe48298083a20100000000,
104'h0839a4bf73427ac58400000001,
104'h663b6d057621dcc14300000000,
104'h0412c701252250454400000000,
104'h66d07b20a0518019a300000000,
104'h54dc0840b8dca784b900000000,
104'h00b5ec886b384da770ee3a2fdb,
104'h00ac914c59db87deb788192b10,
104'h348f51ea1ed5db26abffffffff,
104'h6685d5ae0bb294726500000000,
104'h90fab4b0f59e30123c6484a2c9,
104'h2c2f1fb35e0a28191400000000,
104'h60420307840941ab1200000000,
104'hbc67dc67cfc2316e8400000000,
104'h04713bdbe2902ee62000000000,
104'h34bca7967928ced151ffffffff,
104'h34fd5ad6fa543c85a8ffffffff,
104'h340b17cb16e0aa5ac100000000,
104'h30e80468d06b9103d700000000,
104'hbc804a5200d315e8a600000000,
104'h9c0bf1bb178fb0981f0bb09817,
104'h9c9e2f3a3c49e7179308271210,
104'h00fe1cb8fca9b94253a7d5fb4f,
104'h6693954a270d133f1a00000000,
104'h04afac105f785ec1f000000000,
104'h60f2f614e5200b814000000000,
104'h66bc9f2c794ba68d9700000000,
104'h669401de287ad8b5f500000000,
104'h00133a39269263e024a59e194a,
104'h602bebb957daf778b500000000,
104'hb8603223c0b573bc6a00000000,
104'h66e8756cd087f4280f00000000,
104'h006b9897d77cb8d9f9e85171d0,
104'h6019bb8933a7c6e04f00000000,
104'h665287fda5f9d7b2f300000000,
104'hb8b6c1566d7eef7dfd00000000,
104'hbc498f8593b4b2866900000000,
104'h9c48bce391b851967008108210,
104'h0453df19a795a5502b00000000,
104'h348922fa1290d08e21ffffffff,
104'h661b336736c981cc9300000000,
104'hb8be73287c82ab7c0500000000,
104'h00d481d8a99b4b74366fcd4cdf,
104'h60a3c3ba47cc99409900000000,
104'h54dd649cbaffb388ff00000000,
104'h2c670dbbcef0a472e100000000,
104'h047e469bfc4e55019c00000000,
104'h080a38f51406c7710d00000000,
104'h66fd4f84fa64b09bc900000000,
104'h9032e7f7657f4857fe4dafa09b,
104'h04ee0fc0dc2ee8d35d00000000,
104'h3435040b6ab0d5006100000000,
104'h3469ec7fd3523de5a400000000,
104'h08e4093cc84e5f099c00000001,
104'h949d4baa3a7549cdea00000000,
104'h0077125beea0b7ce4117ca2a2f,
104'h00d57fecaa61fc47c3377c346d,
104'h288ba4ee171fec6b3f00000000,
104'h08fb74b4f6fd56cefa00000001,
104'h54133d4526c861bc9000000000,
104'hbc271a2f4ed0e89ea100000000,
104'h34b79a6a6f47b05d8fffffffff,
104'h94b791446fa20ab64400000000,
104'h2801ca2d03dd40a8ba00000000,
104'h281c17a33852dbcfa500000000,
104'h084ff5139f8aa6bc1500000000,
104'h2c39b3b57308fc651100000000,
104'h5465ea6dcbefbe74df00000000,
104'h2819a0a933560ab5ac00000000,
104'h04246c4748ee876add00000000,
104'hbc4c7a6b98dddebabb00000000,
104'h2cb33b6866f2c0fee500000000,
104'h602e29a35cb686306d00000000,
104'h6629e36553794649f200000000,
104'h90f68fc2ed7e0097fc888f5511,
104'h0483468006332a296600000000,
104'h3042f2f185e1bb26c300000000,
104'h9067e9cdcfe09336c1877afb0e,
104'h60842a1c0813ccdb2700000000,
104'h9c1b011336bf57d07e1b011036,
104'h907d88f1fb69f271d3147a8028,
104'h60963ae02c295a135200000000,
104'hb8c08bda81224a654400000000,
104'hb8a04c8040bea3d87d00000000,
104'h04d14404a209d0f31300000000,
104'h046a3dffd43742bd6e00000000,
104'h905f835bbf809c1601df1f4dbe,
104'h9cff7628feb8e41e71b8640870,
104'h34c0c88a8117d78d2fffffffff,
104'h04948688294c31179800000000,
104'h9496eafe2dc580d08b00000000,
104'h2c80b76c01cdea849b00000000,
104'h604f86e39f69e31dd300000000,
104'h006e53dfdc77c501efe618e1cb,
104'h34e82924d022d36f45ffffffff,
104'h340db5ab1bdd04e8ba00000000,
104'hb8233b6f46a8ac845100000000,
104'h2c57115faef6da58ed00000000,
104'h6019b02f33b10ad66200000000,
104'h342702454e9c7d2c3800000000,
104'h94d56e8eaa1348a32600000000,
104'hb8c1d668838308fe0600000000,
104'h54607e7bc02ab9e55500000000,
104'h9c899a9813a1192e4281180802,
104'h0474f4a1e9b2a8566500000000,
104'h90f2e65ee59224d42460c28ac1,
104'hbcb99e6a73180f793000000000,
104'hbc84680808559ad1ab00000000,
104'h9c376e056efd1882fa3508006a,
104'h546d309fda85bdba0b00000000,
104'h5473a65de76a5675d400000000,
104'h2cfdbff2fbe23ff0c400000000,
104'hb85ac71db5e9c206d300000000,
104'h600fd08b1fca9f8e9500000000,
104'h28e838b2d08775b60e00000000,
104'hb828e3b75104426f0800000000,
104'h9036b8496d7429c1e842918885,
104'h54e38d82c7e85230d000000000,
104'h946583cbcbc570208a00000000,
104'h00eb80b8d7d5582eaac0d8e781,
104'h2c7e45e7fc8fb0921f00000000,
104'h08985ae4308099820100000000,
104'h3447c2078f55e491ab00000000,
104'h28f33052e683330a0600000000,
104'h90b14058628b135a163a530274,
104'h08b2d810653ef5657d00000001,
104'h2c42b9c585a18de84300000000,
104'hbc7af7e9f5f700e8ee00000000,
104'h08bdc3fc7be3eafac700000001,
104'hbc69d069d3b821b47000000000,
104'h2cdb3d66b613c3092700000000,
104'h08c0c8da816ceba3d900000001,
104'h08d1b932a38a2c501400000000,
104'h0833bb4b673996537300000001,
104'hb810ab4d2155f6cfab00000000,
104'h302b008756fb991ef700000000,
104'h345c545db893a83c2700000000,
104'hbc043c19088907201200000000,
104'h2c366dd36cfb381af600000000,
104'h081de84f3b0bab371700000000,
104'h903f95db7f5f8ba1bf601e7ac0,
104'h6639a2337393e3fe2700000000,
104'h34fd7b5efa9bb1ce37ffffffff,
104'hbc81359002bf3fd07e00000000,
104'h5431ca0b6329df5d5300000000,
104'h303a68f7740ed8cb1d00000000,
104'h9cadd64a5b602ac9c020024840,
104'h2cf589aeeb4970c79200000000,
104'h344f094d9e0f084f1e00000000,
104'h28c2b7c485054d650a00000000,
104'h04900cfc20fd85eafb00000000,
104'h08b9f2067335d3ff6b00000001,
104'h2cdab802b57f4759fe00000000,
104'hbce1e1fec358e5afb100000000,
104'h9c86b9d00d2042134000001000,
104'h284167fb829ffb523f00000000,
104'hbc31068d622239594400000000,
104'h90a7e7024f3101876296e6852d,
104'h94d80326b047fa238f00000000,
104'h9c7850e9f05af4a9b55850a9b0,
104'h30e87148d02a572f5400000000,
104'h3482f232055a3ccfb4ffffffff,
104'h30271b614e12e4fb2500000000,
104'h04b9fe307308c9db1100000000,
104'h60234099461875bf3000000000,
104'h904cdaef9995ef662bd93589b2,
104'h949dc0dc3bf95576f200000000,
104'h28762d37ec2200cf4400000000,
104'hbc1108db22ef45e2de00000000,
104'h3008a49511d9ad2cb300000000,
104'h3045bdfd8b793a7df200000000,
104'h948687540ded1b5eda00000000,
104'h08a02a6e40d6d47ead00000001,
104'hbc4ffe859f7ec601fd00000000,
104'h2892691e24b19ee86300000000,
104'h2c3421ef6866176fcc00000000,
104'h285f51b7be300a736000000000,
104'h6670c421e161c5c5c300000000,
104'h2c1a24a5346e299bdc00000000,
104'h9cecfe64d915eedf2b04ee4409,
104'h548ef7121d182c9d3000000000,
104'h003a7cc774f1f458e32c712057,
104'h607fdeedffa29d744500000000,
104'h08a98a1453da178cb400000001,
104'h0062dee1c55c5bdfb8bf3ac17d,
104'h087bdbd9f730d59b6100000000,
104'h048c925819565955ac00000000,
104'h34021e61049c035a3800000000,
104'hbc739981e7dd1516ba00000000,
104'hbc3040b760a1a96a4300000000,
104'hb878c547f1ffd81cff00000000,
104'h34f480a6e9f8a026f1ffffffff,
104'h66600355c061b125c300000000,
104'h605d36bfba28ebab5100000000,
104'h9c660a19cc5030aba040000980,
104'h60596249b2d7d7d2af00000000,
104'h549ec4bc3ddbe4eab700000000,
104'h949ff5503fdbd43ab700000000,
104'h08087f2d106e95e1dd00000001,
104'h6609e0a513f4103ce800000000,
104'hbc7fd217ff1b41493600000000,
104'hbc6adfcfd5bfd6f87f00000000,
104'h00804ee400a3d69e4724258247,
104'h60b5051c6a51ab47a300000000,
104'h085debc5bbf0b31ce100000000,
104'h08f30598e67a23c5f400000001,
104'h04632f9fc675ddc1eb00000000,
104'h3065450fcaa686ce4d00000000,
104'h90001e2500c2034884c21d6d84,
104'h9ccda20a9bef2680decd22009a,
104'h30f5e3bceb33322d6600000000,
104'h54b601da6cb17cb66200000000,
104'h002b4197568d56aa1ab8984170,
104'h003d9c8b7bd2070ca40fa3981f,
104'h0495b99c2bee76bedc00000000,
104'h30b908e47281e2dc0300000000,
104'h66637a7dc65cae23b900000000,
104'h9c310875622429474820084540,
104'hbc520ba1a4e9ea56d300000000,
104'h2c8c138618af0b225e00000000,
104'h9cddb936bb2966955209201412,
104'h34eea528dda4ad0e49ffffffff,
104'h28b5c0286b72e7d7e500000000,
104'h2c9e47243c7fc367ff00000000,
104'h66a13a22422fb8db5f00000000,
104'h54735e09e62fee475f00000000,
104'h60c0c990812d661d5a00000000,
104'h08a5b51e4b01d58b0300000001,
104'h94d905a0b2b239d86400000000,
104'h947fca75ff0f04cf1e00000000,
104'h9411a63f23cf780a9e00000000,
104'h9c44dad38911876d2300824101,
104'h60557013aa2d5a6f5a00000000,
104'h3055adc9ab3744856e00000000,
104'h043ee08d7d4ccc7f9900000000,
104'h2c6021a3c0511aefa200000000,
104'h343d99d97bfae77af500000000,
104'h5425776b4a79bd49f300000000,
104'h30608ee1c1722e5be400000000,
104'h28235eed46104def2000000000,
104'hbcf0ef50e16589dfcb00000000,
104'h662bc2b757a2bafc4500000000,
104'h90c9d39693f1047ee238d7e871,
104'h28b754126e23da4f4700000000,
104'h9418a8db312c46795800000000,
104'h347ed70dfd8945801200000000,
104'h94f25d0ee4dad1c8b500000000,
104'h90a72e724eacf5ec590bdb9e17,
104'h90e94adad275fe29eb9cb4f339,
104'h948c27ce180ea0b31d00000000,
104'hbc8fe5aa1f8cb5181900000000,
104'h54f6076eecd0d2aaa100000000,
104'h9c9425aa2834edd16914258028,
104'h9c45d45d8b0dcc731b05c4510b,
104'h08dfb3c8bf0ae9511500000001,
104'h94e46464c8601e67c000000000,
104'hb8e8d5aed1fa2e50f400000000,
104'hbc002815003b04a37600000000,
104'h902019cb40cc454e98ec5c85d8,
104'h9c65b6b7cb6e8303dd648203c9,
104'h5426c3474d3934877200000000,
104'h30ff1a56fef34122e600000000,
104'h3439f60f73f5bbf4eb00000000,
104'hb845dbc38bda265cb400000000,
104'h30fea2d0fdfb5154f600000000,
104'h00b3ce8467fbb5d0f7af84555e,
104'h289a32f63405dc210b00000000,
104'h60fe9ce8fdc32a568600000000,
104'h60c3f4ac870331990600000000,
104'h04aa13fc5431528d6200000000,
104'h283b46e176f050b4e000000000,
104'h083d2f8d7af32ccee600000000,
104'h04ce853c9d605e33c000000000,
104'h0425e6214b2843395000000000,
104'h60deb42ebda960905200000000,
104'h0417b5092f34c7a76900000000,
104'h9c0bece11772bc07e502ac0105,
104'h2870ec51e1bb6fb47600000000,
104'h3476893fed216e914200000000,
104'h90f2bac0e59b10bc3669aa7cd3,
104'h00c10ff6825e0befbc1f1be63e,
104'hbcd7f9eaaf8bfbde1700000000,
104'h28bee0727db0799a6000000000,
104'h6016ba152db919f27200000000,
104'h667b9edff7ed6aceda00000000,
104'h00588e4fb170c797e1c955e792,
104'h9c0760290ef19c8ae301000802,
104'h34f59862ebc9712692ffffffff,
104'h543395fd67e6d186cd00000000,
104'h54fe54defcd5eebeab00000000,
104'h542cbac3590e8e411d00000000,
104'h9020270d40c5a03a8be58737cb,
104'h289cbdaa39ce94f49d00000000,
104'hbcf0a4f8e10c49351800000000,
104'h30c22e9e847b219ff600000000,
104'h66eba370d76dad0ddb00000000,
104'h90a82a4c501ae5fb35b2cfb765,
104'h043001ff6088eada1100000000,
104'h286b061fd620c5834100000000,
104'h30c736f08e3f997f7f00000000,
104'h3035bc436bd75176ae00000000,
104'hbc039b510714a3912900000000,
104'h046417a1c8fa04cef400000000,
104'h004176eb825ee36fbda05a5b3f,
104'h60f59feaebb840487000000000,
104'h2816cc4d2deb7f34d600000000,
104'h083d45877a1e06613c00000000,
104'hb8bde4c07b6c04bfd800000000,
104'h9c79cda5f39e77523c18450030,
104'hb8469c538dcc45a69800000000,
104'h2cc2fe30853c0d1b7800000000,
104'h30da6dd0b44bf34d9700000000,
104'h2c7789d3ef8a97741500000000,
104'h081f3ec53ef7fac8ef00000000,
104'hb817bbfb2f86f7dc0d00000000,
104'h2c84eb7a09dfa0fabf00000000,
104'h0438e4d571009d8d0100000000,
104'h0809930113215e7b4200000001,
104'h2cfd854afb10c1852100000000,
104'h04c0a32281ab7ba65600000000,
104'h343e3b097cdb627cb600000000,
104'h0428a469514c6c9b9800000000,
104'h904f6c7b9e9600f22cd96c89b2,
104'h001bc623376eed33dd8ab35714,
104'h300fb4cf1f901b222000000000,
104'h9ce72a5cce9ddd083b8508080a,
104'h04ab0ff056b969087200000000,
104'h34d4f1dea9abdb7c57ffffffff,
104'h943ec6897de1d85ec300000000,
104'h5435083b6a1aa3a73500000000,
104'h344a1a0994af48a45e00000000,
104'h28b0afb6611e28673c00000000,
104'h0097b0962f0507150a9cb7ab39,
104'hb874cd63e9577055ae00000000,
104'hb80bc12317590aa9b200000000,
104'h907ef509fd2331cf465dc4c6bb,
104'h6082ff560532f01f6500000000,
104'h0019353732182ef13031642862,
104'h2cae47a05cd0b5f2a100000000,
104'h0450a337a11151972200000000,
104'h28970b2a2ead38605a00000000,
104'h2cf2a714e5df875abf00000000,
104'hb8387be170646d65c800000000,
104'hbc5d079fba7f5d9dfe00000000,
104'h9c597871b23160bb6211603122,
104'h602cb65f596e5d75dc00000000,
104'h609338442601efdf0300000000,
104'h34975ba22e7c27c3f8ffffffff,
104'h0430b78961dc460ab800000000,
104'h00fba274f733511f662ef3945d,
104'h9452e32ba512183d2400000000,
104'h54f444a0e8b5fde66b00000000,
104'h308584d40b7da133fb00000000,
104'h00f9d6b4f3aa3e3654a414eb47,
104'h04b0eef461c45d648800000000,
104'h285f53fbbe9229ea2400000000,
104'h9c1468b5285b8711b710001120,
104'h54356a7f6aabbc9c5700000000,
104'h9cb55a006aca52329480520000,
104'h3060870fc13471ad6800000000,
104'hb86f3787de65e885cb00000000,
104'h60eda134dbaca0325900000000,
104'h34902eb02083258606ffffffff,
104'hb871c73fe376970fed00000000,
104'h08ae91aa5dda1270b400000001,
104'h90006a3500ed78d8daed12edda,
104'h94230363469722422e00000000,
104'h280469e908cfd7ee9f00000000,
104'h54536383a6562db5ac00000000,
104'h5407e0e10f9a126c3400000000,
104'h08ba7a7874032f450600000001,
104'h0836b06d6d2c6e2d5800000000,
104'h3458656fb05cbf2fb900000000,
104'h3427cc994fd8f4ceb100000000,
104'h9cf7c250ef944f6e2894424028,
104'h0439482f72b50fac6a00000000,
104'hbc739bcde74827c19000000000,
104'h9c8b20ba16cae3e0958a20a014,
104'h28ea154cd4d3219ea600000000,
104'h9064ca89c9866e480ce2a4c1c5,
104'h6687d6fe0fae24485c00000000,
104'h54917ca6227a5f83f400000000,
104'h905839cbb05f60b7be07597c0e,
104'h2cff3cdefe58b7e7b100000000,
104'hbc4633638c334da96600000000,
104'h9cacabbe59bb239276a8239250,
104'h543a022d74bb63967600000000,
104'h04b19090631716612e00000000,
104'h2cff9958ffce98be9d00000000,
104'h9cee2560dcf9a7f0f3e82560d0,
104'h6661ccd3c3879d1c0f00000000,
104'hb8ad22fc5a672f9dce00000000,
104'h04a63d424c7cd66bf900000000,
104'hbc448cef89faa07ef500000000,
104'h54560419ac2e1c295c00000000,
104'h30813d840220a5754100000000,
104'hb8ff1f80fe64338fc800000000,
104'h086931c9d28a7d1c1400000000,
104'h945a9e65b5fe0b9cfc00000000,
104'h34a0958641b495ce69ffffffff,
104'h30038c710767b90bcf00000000,
104'h007d8f4dfb1ce9a9399a78f734,
104'hb8aa9e1055b732566e00000000,
104'h2c96cc642d851a840a00000000,
104'h2c729c73e52acbbd5500000000,
104'h3058ccdbb15c4e03b800000000,
104'h28e19182c38573380a00000000,
104'h66edef7cdb2cc97d5900000000,
104'h2892b3e82584ac860900000000,
104'h66853dd40aa94e0c5200000000,
104'h309513162a6c4d21d800000000,
104'h90c3f83087b634906c75cca0eb,
104'h542303334663f847c700000000,
104'hb8ede198db8a49a41400000000,
104'h281e492d3c225af14400000000,
104'h08104bdf20c369a68600000000,
104'h667d06affa2227dd4400000000,
104'h003be389770adcad1546c0368c,
104'h54936626265cd389b900000000,
104'hbc993be632a572984a00000000,
104'h34e606becc47102d8effffffff,
104'h90e41b04c80b5f0516ef4401de,
104'h28f12862e28b09c41600000000,
104'h949985ac3363d54dc700000000,
104'h601097c121bc62107800000000,
104'h08e48b6ac980648a0000000000,
104'h54745a43e801ec8b0300000000,
104'h9415d28b2bb4139c6800000000,
104'hb8ce1a149c712a6de200000000,
104'h2c31e41b63a23d1e4400000000,
104'hbc235225469786b62f00000000,
104'h28e237e4c4e12b6cc200000000,
104'h54f03a1ce06d5221da00000000,
104'h28d50076aa0c74a31800000000,
104'h9087726a0eae7f285c290d4252,
104'h9c57b71bafa3169c4603161806,
104'h305a7039b4551e0baa00000000,
104'h54b867dc70cd52f69a00000000,
104'h6096a9722db198c26300000000,
104'hb8b9bd8a73e64b0acc00000000,
104'h284380c7875caf0db900000000,
104'hb825cdaf4b655bf9ca00000000,
104'h60ccf19e99ff3262fe00000000,
104'h944ba49797833a980600000000,
104'h90a6fc264dab8204570d7e221a,
104'h2cf3914ce7b6cf886d00000000,
104'h9c75d14deb44c6eb8944c04989,
104'hbc16319d2ce5d324cb00000000,
104'h34e6bebacd2fefd35fffffffff,
104'h66623e15c4e52988ca00000000,
104'h2c25dadf4b4a6d399400000000,
104'h045d15ffbaa4fe904900000000,
104'h309c70e238e2ad58c500000000,
104'hb8aa0b665424a1d94900000000,
104'h04642cb3c82e582f5c00000000,
104'hbcc46f1a880a22bb1400000000,
104'h049b06fc367a4b77f400000000,
104'h94385ca57079ac57f300000000,
104'hbc83f12a071056ad2000000000,
104'h302646534c88a1841100000000,
104'h9c20416b408eb70a1d00010a00,
104'h909d412e3a6878e3d0f539cdea,
104'h9caddea45b2d538f5a2d52845a,
104'h28181105302558cd4a00000000,
104'h60362c8b6c2cb8f75900000000,
104'h0428f4615194735e2800000000,
104'hbc19b783336ad5bbd500000000,
104'h0020309140ce22749cee5305dc,
104'h3044a0bd89d97618b200000000,
104'h28395da1724fc3ab9f00000000,
104'h9477ca23ef52800da500000000,
104'h609b725a36a1545a4200000000,
104'h9cd2c262a505ef510b00c24001,
104'h3437904b6f1acda53500000000,
104'h348a70e6147d9165fbffffffff,
104'h34528fbda52540614a00000000,
104'hbc7881ddf1f28182e500000000,
104'h28454bbf8a13b12d2700000000,
104'h94ef922edf7064a5e000000000,
104'h2cbfae1a7f6fb465df00000000,
104'h66001b89000265890400000000,
104'h049a7b5e3455ca25ab00000000,
104'h9c1a205734e5f0aacb00200200,
104'h3403ded5073d7a497a00000000,
104'h2cb797c66f7f3047fe00000000,
104'h2892b68a2549306d9200000000,
104'h007b99c5f78b48581606e21e0d,
104'h2c8c9f4819f9d7eaf300000000,
104'hbcf24af8e4cc529c9800000000,
104'h006ac09fd5e237e2c44cf88299,
104'h94dd88d2bb2b1a8d5600000000,
104'h346958d9d2b60f2c6c00000000,
104'h66ba557e740a99691500000000,
104'h9cae09005cd0f066a180000000,
104'h94eb03e6d64932299200000000,
104'h5450e0e3a110dded2100000000,
104'h54b223b6642bad8d5700000000,
104'h28542b0da8a0a5da4100000000,
104'h04ea2d5cd42df60d5b00000000,
104'h5456f8c9ad0dfe0d1b00000000,
104'h6625ee014b7593e7eb00000000,
104'hb88e6e221cc7601e8e00000000,
104'h00a5b3944b61e917c3079cac0e,
104'hbc51cde9a3dda56abb00000000,
104'h044d38c19a762d57ec00000000,
104'h344545a58aa563104a00000000,
104'h308650f00c992a263200000000,
104'h90ef79a4de9405e8287b7c4cf6,
104'h28bc54507866b6bfcd00000000,
104'h3445d0f38b74ae91e900000000,
104'h08dc4bceb80ef41f1d00000001,
104'h9c7b815bf7d0cd64a1508140a1,
104'hbc05dd150bff48fefe00000000,
104'h601f5b6b3e287e815000000000,
104'h9058f691b1511ddda209eb4c13,
104'h9454566da856a5c1ad00000000,
104'h908c3b6c18ba58f4743663986c,
104'h34b0dc6c613ccac179ffffffff,
104'h30b82f94707b9a43f700000000,
104'h3010d6392192b4da2500000000,
104'hb88323b6068837821000000000,
104'h3466775bcc75c72feb00000000,
104'hb899e13c33e3f82ec700000000,
104'h2855ca1fab141c952800000000,
104'h6621165342f29186e500000000,
104'h6026fb934d8f63aa1e00000000,
104'h088b81e61734e2836900000001,
104'h945b6783b6f37acce600000000,
104'h9000dfa301afefe05faf30435e,
104'h00f16476e2dccc16b9ce308d9b,
104'h2c4193f583f9a01ef300000000,
104'h3022cfbf452a69655400000000,
104'h66b3180666a737744e00000000,
104'h662a596754d7e852af00000000,
104'hb80125c5029993de3300000000,
104'h305b9037b7dafe3ab500000000,
104'h307fa3ddff63291dc600000000,
104'h2c99adc033a0dc3c4100000000,
104'hbc3951b972c3bca88700000000,
104'h08f9224af2874b300e00000000,
104'h94573385aef5e1bceb00000000,
104'h6617e0e52f6d87b5db00000000,
104'h284cbe2f994a35599400000000,
104'h08786b59f038de257100000000,
104'h08f4c362e94c5a359800000001,
104'h04eb9e34d7e9069cd200000000,
104'hb88b1d88166db4cfdb00000000,
104'h9cd53cc2aa9840f8309000c020,
104'h042f1bd15ef1e762e300000000,
104'h34d73d0eae8330d206ffffffff,
104'h045aae25b5990dec3200000000,
104'h662fd3e75ff4798ae800000000,
104'h087a5133f443ba298700000000,
104'h54d640d4acb01a386000000000,
104'h9091ba64238caf90191d15f43a,
104'h30225a27443a89bd7500000000,
104'hbc9943e832145f652800000000,
104'h308ad8e6151792af2f00000000,
104'h940018a700fa249cf400000000,
104'h28c664e08cdcef6cb900000000,
104'h607f2051febf3ff67e00000000,
104'h665b60a3b6b4a6126900000000,
104'h2c28ab4d518f93ee1f00000000,
104'h9c6a7577d4ab247c562a247454,
104'h2860decbc1ac20c05800000000,
104'h303fdf697fe51c44ca00000000,
104'h2c2ae0b755734069e600000000,
104'h28f77946ee991eca3200000000,
104'hbcf6c3b8ed42a2a38500000000,
104'h083f889b7f68f927d100000001,
104'h00dc3340b82f08eb5e0b3c2c16,
104'hbc0649b10c76d039ed00000000,
104'h60eddf7adb4dc27b9b00000000,
104'hb89e3b963c51fc99a300000000,
104'h3411a951230be8531700000000,
104'h94a52c184a97a6a42f00000000,
104'hbc898e6e13cf592a9e00000000,
104'h90ba03be74e32278c65921c6b2,
104'h2c19554132dd7580ba00000000,
104'h08cd51d89a6a0bf1d400000001,
104'h0874f8f5e9439b918700000000,
104'h08989872316022a7c000000001,
104'h0863d577c73d63577a00000000,
104'h2c88585410fee5fafd00000000,
104'h2cc4936e89549a8da900000000,
104'h2c24dd1149ccf1049900000000,
104'h545dd44fbb3700b36e00000000,
104'h90c5c8ec8b8116a40244de4889,
104'h94279e3d4ffdc302fb00000000,
104'hbc1c60f9389d3d723a00000000,
104'h94798829f362b877c500000000,
104'h00e098fec19cfbcc397d94cafa,
104'h0449a5bd931f5dcd3e00000000,
104'h9cacdf8c5953f3cfa700d38c01,
104'h60683367d0719181e300000000,
104'h94d4a9eca9d7ef54af00000000,
104'h90640251c8820fce04e60d9fcc,
104'h04c1c02a8312bbf92500000000,
104'h0483a4660728aeb35100000000,
104'h2c24491548d7c71aaf00000000,
104'h94ff5856fe4a59e99400000000,
104'h60019635031979d33200000000,
104'h2c67b58bcfccceec9900000000,
104'h086dafd9db9a55003400000000,
104'h66e5182ecadc18f8b800000000,
104'h907ba10bf735cd3d6b4e6c369c,
104'h00bbcd3077fdcd0afbb99a3b72,
104'h60b08396619ce6e43900000000,
104'h3440fe3b812e05e15c00000000,
104'h04054c0b0a2292154500000000,
104'h902c5dbb58021ff3042e42485c,
104'h604355b186f3c6a8e700000000,
104'h66f292dae58d357e1a00000000,
104'h6047ae958fd7603aae00000000,
104'h6694658628825a800400000000,
104'h2c792385f251ba2ba300000000,
104'hbc0eaa6d1dd098b2a100000000,
104'h9c7d0c0bfac80b909048080090,
104'h2856eef7adb4ab946900000000,
104'h9cf6d674edff834cfff68244ed,
104'h5490e55021fc7c5ef800000000,
104'h28de53cabc1423f72800000000,
104'h94e89068d1f85e10f000000000,
104'hbcb8c3de71c35fec8600000000,
104'hbc3d2fe97a560963ac00000000,
104'h04c0a13681a6754a4c00000000,
104'h0488ec3e11e158d2c200000000,
104'h30c82d2290b889ea7100000000,
104'h28b1429462e6c49ccd00000000,
104'h9062bbafc544876d89263cc24c,
104'h342c30d758b39ebc6700000000,
104'h08a0bfa44116b72b2d00000001,
104'h54a621b24c700eefe000000000,
104'h286a9691d58e1e3e1c00000000,
104'h28949892294ecead9d00000000,
104'h344614bf8ce99986d300000000,
104'h08619da5c3cea5369d00000000,
104'h0412d13d25ecb9a0d900000000,
104'h349be9d03789a38413ffffffff,
104'h900931d512b85ee470b16f3162,
104'h9057d2c9afce20569c99f29f33,
104'h6008371510731571e600000000,
104'h60acf6f259fd7424fa00000000,
104'hbcfe0846fc1d311f3a00000000,
104'hb8fca97ef96c752dd800000000,
104'h08f73f76eeaca98e5900000000,
104'h906d1e59da41b36b832cad3259,
104'h3420f573414cb61b9900000000,
104'h66c556288a8d74981a00000000,
104'h60c98dc4935d29ddba00000000,
104'h0095ca5e2b9770362e2d3a9459,
104'h902c42bb588d8fb21ba1cd0943,
104'h2859d927b31e4b7d3c00000000,
104'h0893715e2630063b6000000001,
104'h90fdf16afb04d56b09f92401f2,
104'hb81da57d3b9fdbcc3f00000000,
104'h04f67ed6eca902b85200000000,
104'h083165a36257ea87af00000001,
104'h94d395d6a7e0a9e4c100000000,
104'h2c6bbf1bd714b4432900000000,
104'h30fd5f98fa57ff2baf00000000,
104'hb89591f02b1e3ea13c00000000,
104'h040546090acdd0869b00000000,
104'h2ceb9cf2d795aefa2b00000000,
104'h94b7dfce6f6981b5d300000000,
104'hbcc549aa8a62a66bc500000000,
104'h04db9c5cb726c82f4d00000000,
104'h2c663867cc1c5dcf3800000000,
104'h60482fd9901327352600000000,
104'h94868c2e0d0a81c31500000000,
104'h2cc2bf3285d92bbeb200000000,
104'h08ddf6d4bb19cea53300000001,
104'h28cacc1495d5688aaa00000000,
104'h34bd84de7b606c8bc0ffffffff,
104'h0843e0ed87b132166200000000,
104'h9c84299c088e0b561c84091408,
104'h30a7fce44f3f1a9b7e00000000,
104'h947a0b1bf463bea3c700000000,
104'h042ebfe95d152e132a00000000,
104'h9c5e8e23bd0f99cb1f0e88031d,
104'hbc1556a72a20ee3f4100000000,
104'h04b522406a080be91000000000,
104'h34f32688e6310e9962ffffffff,
104'h549ccdc039c2fbda8500000000,
104'h34c739ba8e30f05b61ffffffff,
104'h2cbe79b07c64a43dc900000000,
104'h542a6b2b5491de842300000000,
104'h909dfdda3b422f6b84dfd2b1bf,
104'h66d25282a41e09cf3c00000000,
104'h9059eccdb3d41380a88dff4d1b,
104'h0450f031a13144b76200000000,
104'hb8a61fd04c742e5be800000000,
104'h9cbd195e7a137f792611195822,
104'hbc8d02f21a03a1950700000000,
104'h04afa3f85ff10410e200000000,
104'h9c43a10187546e89a840200180,
104'h04c152ac82ac723a5800000000,
104'hbc1c6f8538f2d256e500000000,
104'h607580e5eb867b700c00000000,
104'h2c64dacdc9aa61d65400000000,
104'h543d8ecd7b575ef3ae00000000,
104'h00b991e273e2e5a6c59c778938,
104'h00010d5302d625b8acd7330bae,
104'h281d92933bb0f6226100000000,
104'h9056aa21ad299e81537f34a0fe,
104'h04dff56abf3657676c00000000,
104'h3059dba5b3bf19c67e00000000,
104'h9c1c79b538ae154e5c0c110418,
104'hbcc94d089222e5c74500000000,
104'h2862d17dc5405f778000000000,
104'h54da0a38b4568a7dad00000000,
104'h28d0ad90a17a2539f400000000,
104'h34eb6be2d6e0c5a4c1ffffffff,
104'h00aa897a550471b508aefb2f5d,
104'hb807c3710f9346ba2600000000,
104'h663f37897ef787c2ef00000000,
104'h54ddc710bbc22af88400000000,
104'h30a22cc444e5be00cb00000000,
104'hb89ebdaa3d69395dd200000000,
104'h00888cfa117a1acbf402a7c605,
104'h60ed6af0da7adea5f500000000,
104'h3054f6b7a946b03d8d00000000,
104'h2cc9bb489354e949a900000000,
104'h541e0f473c1eb8333d00000000,
104'h00252fe34a1705872e3c356a78,
104'h083bceb7771870493000000000,
104'h088c0aa81856f95bad00000001,
104'h08a78bd04f12b5d92500000001,
104'h900f3a491e6ea07fdd619a36c3,
104'h663ac821755a6203b400000000,
104'hb85b062db65fa873bf00000000,
104'h3498bbf231cb659e96ffffffff,
104'h08a67a824c090c711200000001,
104'h344ea2559d89a54a1300000000,
104'h66e79434cf2a51735400000000,
104'h9c76c511ed2d95635b24850149,
104'h60782ceff0708237e100000000,
104'h30ea48b4d40096030100000000,
104'h2817a71d2f88eb381100000000,
104'hb8cdb88a9ba50f064a00000000,
104'h90f559eceaf596b4eb00cf5801,
104'h9c0452a108464c0b8c04400108,
104'h082fbd4b5f1f88a73f00000000,
104'h66d613beac2c18695800000000,
104'h60f455dee8e2bacac500000000,
104'h28d48374a94e1b419c00000000,
104'h542c6119588fd89a1f00000000,
104'h66ca400e9442f36b8500000000,
104'h66624125c41fbb573f00000000,
104'hbc414a9782a713844e00000000,
104'h2c4ba8ed9714a5f72900000000,
104'h34ec12d8d8d75deaaeffffffff,
104'h9024881d4945413b8a61c926c3,
104'h2cfd4362fa9b80b83700000000,
104'hbcc6b7228d8d579a1a00000000,
104'h343a4d7f741c11cb3800000000,
104'h602a6327542051554000000000,
104'hb854b539a9406abd8000000000,
104'h28bb3a1a76f97064f200000000,
104'h34d61d5eac5044e9a0ffffffff,
104'h00ae56a65ca5cc844b54232aa7,
104'h2cab137a5675156fea00000000,
104'h0044ec3789640f35c8a8fb6d51,
104'h9c189bdb31772927ee10090320,
104'h28a7b2f64f55efadab00000000,
104'h94a87d8850d280aea500000000,
104'h34c713d48e3f6eed7effffffff,
104'h34584e51b0ff6c62fe00000000,
104'hb86c147bd80fd3ad1f00000000,
104'h00173ec12e8ae85e15a2271f43,
104'h66660357cc30666b6000000000,
104'h345ea623bd5ab87fb500000000,
104'h6680e3920154ed63a900000000,
104'h54714e83e239445f7200000000,
104'h08b0991a6149e8919300000001,
104'h008d80ae1b8533580a12b40625,
104'h089cd49c39fc8db0f900000001,
104'h081dd0313ba0c88c4100000000,
104'h6679bf83f3b8843c7100000000,
104'h30b4a754697cfed3f900000000,
104'h00d967f8b2576175ae30c96e60,
104'h005e9329bd5c64c9b8baf7f375,
104'h94e1ececc3dde450bb00000000,
104'h08974f782ea9b8ca5300000001,
104'h08146a0928c2f18e8500000000,
104'h34ed92ccdb7e44f5fcffffffff,
104'h9090a3ba21dc4facb84cec1699,
104'h30219a754333fb236700000000,
104'h2c81732c02ad22e25a00000000,
104'hb84a767d941f50f13e00000000,
104'h001df24b3b92292c24b01b775f,
104'h044e15ad9c4cdbb99900000000,
104'h346b67c3d607b64b0f00000000,
104'h66b8119670deac9abd00000000,
104'hb8abf2fe57056fb70a00000000,
104'h34bb3a8076656c6fcaffffffff,
104'h3025f82b4b2bc8ab5700000000,
104'h08e9e37ad35137d3a200000001,
104'h04b04c34603f3e277e00000000,
104'h66f0ee4ee1563b23ac00000000,
104'hbc2f20c95e2d52e35a00000000,
104'h9c61978bc3610e7bc261060bc2,
104'hbcedb04edb974b5c2e00000000,
104'h2c560279ac76d1b7ed00000000,
104'h0080a9f6019ea9d03d1f53c63e,
104'h347c8525f99d08703a00000000,
104'h909d5daa3a6f6a3bdef23791e4,
104'h08d5b45caba536084a00000000,
104'hb811a81923c3fe568700000000,
104'h60312fab62783997f000000000,
104'h00c89eaa915f099fbe27a84a4f,
104'h9c352d5d6a3d69fb7a3529596a,
104'h0087fb8e0f36dd536dbed8e17c,
104'h947cc67df97971cdf200000000,
104'h34d249aca4ceb46a9dffffffff,
104'h661902d73200eb6b0100000000,
104'h9019d0b733f9afa4f3e07f13c0,
104'h5480a4f8015abcf1b500000000,
104'h343041136003917d0700000000,
104'h08bab62c75ee343adc00000001,
104'h309f1ff03efb3a2ef600000000,
104'h044fd27f9f18e2e33100000000,
104'h2854f33da99ae3b63500000000,
104'h544e34bd9c083a491000000000,
104'h04d32d9ea60a1dd11400000000,
104'h946c8271d9f2e784e500000000,
104'h66c8da86917589f9eb00000000,
104'h041757e72e0def771b00000000,
104'h28c60a208c3857697000000000,
104'h28f5942ceb598ab7b300000000,
104'h0873fd57e7137f212600000000,
104'h082f650f5e21c1a34300000000,
104'h907e11d5fcaebfd85dd0ae0da1,
104'h0884131408cec8569d00000001,
104'h94176e072e5f5a0fbe00000000,
104'h2cfa8d8ef5611aafc200000000,
104'h90c96d1a92f08bfee139e6e473,
104'h34b8b68871b558446affffffff,
104'h9cf6cafcede9cda4d3e0c8a4c1,
104'h904d6ecb9a6be079d7268eb24d,
104'hb83f90557f8eccba1d00000000,
104'hb87961e7f2102e632000000000,
104'h2cb1be94639528c02a00000000,
104'h6642922385dbf4e2b700000000,
104'h9072bbe3e54beef19739551272,
104'h54dea48ebd31fa916300000000,
104'h604d7f2f9ab0d6446100000000,
104'h54bfecf47facb5ca5900000000,
104'h9c517c23a2af3b7a5e01382202,
104'h90d139e2a25ca8adb98d914f1b,
104'h9c6e4f2ddc84dd0e09044d0c08,
104'h54ac60a258927d122400000000,
104'h2cb829767008573d1000000000,
104'h30578941af50e097a100000000,
104'h94c0fcec814d60019a00000000,
104'h9cd53a8aaa4220998440208880,
104'h0032683d64e2c316c5152b5429,
104'h9093260a26cd86309b5ea03abd,
104'h9c9462d028a61dfa4c8400d008,
104'h6683b40e07a8723e5000000000,
104'h54eca8d4d9e95be6d200000000,
104'h346e4fa1dcff395afe00000000,
104'h2ca2e7364565f1d9cb00000000,
104'hbcc2728c8411bfe32300000000,
104'hb8d5a7a0ab39da8f7300000000,
104'h00f97160f2dfd5f2bfd94753b1,
104'hb80bfc8117ea5280d400000000,
104'h34530767a64153678200000000,
104'h90efed00df2853ed50c7beed8f,
104'h2c78a2abf185f3d80b00000000,
104'h307da10dfbd2d2cea500000000,
104'hb8536ffba678f2a9f100000000,
104'h30d34d52a672b8e1e500000000,
104'h902126e1426466efc845400e8a,
104'h668ddf3c1b2ca1a35900000000,
104'h909395aa27705f8be0e3ca21c7,
104'h945e68f7bce4564cc800000000,
104'h0886ed600d79bf15f300000001,
104'h66444d6f880e09df1c00000000,
104'hbc9acdd4353cd7eb7900000000,
104'hb8982c4e30695511d200000000,
104'h28ba118c746fc829df00000000,
104'hbcd38e04a7a1f2604300000000,
104'h945d59d9ba2895a95100000000,
104'h9cc14fba82923a0a24800a0a00,
104'h04145ac528ab0a0a5600000000,
104'h9482cf5c05a35e0a4600000000,
104'h30a1e71a437a4ea9f400000000,
104'h5495d7982b87661c0e00000000,
104'h60b6bc666d4a489d9400000000,
104'h90c74bd88e48ebbb918fa0631f,
104'h90170ef52e2cb4c5593bba3077,
104'h30be944a7d6c9625d900000000,
104'h9cb6d5d26d1603bf2c1601922c,
104'h548dc9d61ba056524000000000,
104'h0818d6cb3195f5e22b00000000,
104'h6072a22fe53463056800000000,
104'h34fc726af85ff74fbfffffffff,
104'hb8b41bb86859f4b3b300000000,
104'h90262ffd4cff3bdcfed91421b2,
104'h3448e9a591e3c19ac700000000,
104'h00cf098c9ed29b2ca5a1a4b943,
104'h54b29fde650439b90800000000,
104'hbc0677e90c2c2c995800000000,
104'hbc399f0f734582c78b00000000,
104'h60133e9b2630a33b6100000000,
104'h9475c0a5ebb734446e00000000,
104'h349ef7f03dd269f0a4ffffffff,
104'h2ccfc2cc9f0dd36b1b00000000,
104'hbc3860f570047f590800000000,
104'h90677471ce300f3960577b48ae,
104'h54786573f00111cb0200000000,
104'h048aa13c156dbc67db00000000,
104'h28d5ebf8ab3fdb657f00000000,
104'h00a8bd9c515c9173b9054f100a,
104'hbcf461d0e8783e01f000000000,
104'h606f52bfde16a2992d00000000,
104'h04f90706f2cb1f3e9600000000,
104'h307b2a8ff6569dd5ad00000000,
104'h5432fa6965f08478e100000000,
104'h60ca3bb494adc6e25b00000000,
104'h042205814404eec90900000000,
104'h90da55a2b4cfb33c9f15e69e2b,
104'h66a8289c5052770da400000000,
104'h28208c7f41afc6225f00000000,
104'h60f1e6c4e331a9e16300000000,
104'h284565398aec6c8cd800000000,
104'h9c6151cbc2de23a2bc40018280,
104'h0851c17ba3c419388800000000,
104'h0087d6340fdaec68b562c29cc4,
104'h54b88bb2719000a42000000000,
104'h34fac752f542941585ffffffff,
104'h04e9230ad28095080100000000,
104'hbc8eab301d1f0e413e00000000,
104'h00d6876ead17c2612fee49cfdc,
104'h304546998aa54e484a00000000,
104'h049f458c3e9cea6c3900000000,
104'h00fa6916f4f0a346e1eb0c5dd5,
104'h004222cf8486a0a60dc8c37591,
104'h309b78f63699d4183300000000,
104'h9c0b8961179626482c02004004,
104'h2c75bf47eb45fb5b8b00000000,
104'hbc27b4314f20a6534100000000,
104'h28e773d0ce0923691200000000,
104'h08859ae80bc2317c8400000001,
104'h547f8923ff38a25f7100000000,
104'h30f69df6ed767a45ec00000000,
104'hbc583887b00936191200000000,
104'h6636f2856dd350e6a600000000,
104'h28384e097014e0332900000000,
104'hbc4ace7f95e0df5ec100000000,
104'h08c734768ea482064900000000,
104'h005c5493b8cba5689727f9fc4f,
104'h30dfc15abf5938b5b200000000,
104'h2c06402b0c6c347fd800000000,
104'hbccdc1029b9179142200000000,
104'h54b751726e60abe1c100000000,
104'h6002427904a5ebc44b00000000,
104'h9c9a79583433f4876712700024,
104'h948aa38815da0920b400000000,
104'h342fc5875fcebd2e9d00000000,
104'h30565cc1ac9c75443800000000,
104'h66820c6a042e36555c00000000,
104'h9c178d6b2f731c0de6130c0926,
104'h28a5592e4a1c8e353900000000,
104'h344a479394af0d145e00000000,
104'h08ea17bed4672ccbce00000001,
104'h60ae9c065dc417b68800000000,
104'h34f100c8e2ceafd29dffffffff,
104'h9c41665182e02712c040261080,
104'h308bc5b617aca6c85900000000,
104'h947fd8bfff1e5e013c00000000,
104'h2c167cb72c0b0ee71600000000,
104'h2881c85a0371f31fe300000000,
104'h9cb5ccb06ba98f2a53a18c2043,
104'h5436b8f16d24ccc94900000000,
104'h9ca5d9564b2c74535824505248,
104'h04d1a90ca385dd1a0b00000000,
104'hbc85ef0e0b716cd7e200000000,
104'h342f9dfd5f233df14600000000,
104'h2c4cef0999c604f48c00000000,
104'h9cc4efcc89ac0ce658840cc408,
104'h28527b2fa47be2a9f700000000,
104'h605d5547ba560757ac00000000,
104'h2898e22e3116c1ad2d00000000,
104'h28baaff67562e661c500000000,
104'h6643cb7387102f812000000000,
104'h08de9828bd217add4200000001,
104'h34e7a328cfed075edaffffffff,
104'h008aa8ea158689680d11325222,
104'h001dc63b3b20ae41413e747c7c,
104'hbc438c07873966617200000000,
104'h94896e5412fa0ee4f400000000,
104'h04e2c60ac5b051e06000000000,
104'h04395de3729655c62c00000000,
104'h3483424006b893c471ffffffff,
104'h90124c1324956d222a8721310e,
104'h28549eb7a98657a80c00000000,
104'h00ae10d05c0c38f518ba49c574,
104'h90a13834422848e7508970d312,
104'h08db90c4b7f092f8e100000001,
104'h3412f64b25faee9ef500000000,
104'h30ab695e56fb06a8f600000000,
104'h0402d7450577c7a9ef00000000,
104'h9cb55cca6aba4d4474b04c4060,
104'h605f3c2dbe7c26a3f800000000,
104'h28027df3045489c5a900000000,
104'h9c74f4cfe9e3cde8c760c4c8c1,
104'h34c81c82903244e964ffffffff,
104'h90a70bb84e134b9726b4402f68,
104'h04df70e8be8f29281e00000000,
104'hbce15234c2ce15889c00000000,
104'h9ca6084c4cac7ec258a4084048,
104'h0451ac4fa374655be800000000,
104'hb8b2f0a0652167b34200000000,
104'h54b41cd46884d4660900000000,
104'h088ca48c1984dbb20900000000,
104'h903d91517bfdb7ccfbc0269d80,
104'h664bb77d976d6443da00000000,
104'hb8f16e10e2fa3c64f400000000,
104'h04d6419cac82989a0500000000,
104'h28edda1edba742cc4e00000000,
104'h04200bdb401c59bb3800000000,
104'h28facb46f56bfb61d700000000,
104'hb89b7be036abce5a5700000000,
104'h5467d217cfe2423cc400000000,
104'h30c7401c8eea1ef8d400000000,
104'h6004a5d909fabb3cf500000000,
104'h2c84bbb80988f1d01100000000,
104'h34c070988068adfdd1ffffffff,
104'h60a332a046e0a6dec100000000,
104'h303bdb257731a1d76300000000,
104'h94cbb58297d853deb000000000,
104'h2859d907b3fcb9eaf900000000,
104'h60b9cdc87303804b0700000000,
104'h349b348a367dd111fbffffffff,
104'h546ce99fd9b1a1626300000000,
104'h2cd0dabea11855e73000000000,
104'hbcbe87f27d6b561fd600000000,
104'h0470e76fe195e6c82b00000000,
104'h3089246e1219633d3200000000,
104'hbc9a7122348cadd21900000000,
104'h044be38197d16f3aa200000000,
104'h5494152a28d17ce0a200000000,
104'hb8f6fe52ed047e510800000000,
104'hb8514393a211a98f2300000000,
104'h604ceed1998b2e7a1600000000,
104'h904a4b239470a937e13ae21475,
104'h94045ba908cbb3789700000000,
104'h28b3256c66c56cf88a00000000,
104'h9496c4442df592c4eb00000000,
104'h00dd02b6bad37daca6b0806360,
104'hb867ecd1cf0f1f991e00000000,
104'h944e96119d9bd7f03700000000,
104'h00b20a3a6450b6f5a102c13005,
104'hb8df2144bea188204300000000,
104'h5462ae2fc509bb911300000000,
104'h08e040e0c0be06587c00000000,
104'h60d47314a80b51eb1600000000,
104'h0022782f44e15274c203caa406,
104'h6011681d2254dc3fa900000000,
104'h34607d3bc0d9d00eb300000000,
104'h280a3d31147e3689fc00000000,
104'hb85d44d3baffe286ff00000000,
104'h30ee2efedc1bb2853700000000,
104'h28c0ce80816148f5c200000000,
104'h048fb2f01f17d3ad2f00000000,
104'h347fb093ffc83a389000000000,
104'h3481e33403becb407dffffffff,
104'h34596413b2ba40ea7400000000,
104'hb85aaab3b5f7b438ef00000000,
104'h28b950cc724ad7699500000000,
104'h6645b11d8be78f52cf00000000,
104'h5406994f0d5dc3cfbb00000000,
104'h9cd406d8a8f9ff0af3d00608a0,
104'h302ea6e35db533f86a00000000,
104'h28b49116690bc39d1700000000,
104'h90f67594ece79980cf11ec1423,
104'h54c135c28232f7056500000000,
104'h665ea033bd1945c73200000000,
104'h948cc784196108ffc200000000,
104'h54262c474c15c5e32b00000000,
104'h305db1cdbbda7b06b400000000,
104'h0438161d7024feb54900000000,
104'h044164c782405c578000000000,
104'h608f9cc21fb808d47000000000,
104'h2ca4815c49a785ee4f00000000,
104'h08df4e04bec9cca09300000000,
104'h089bc53a37f99686f300000001,
104'hbc06d26b0d8f5e341e00000000,
104'h08c9b6cc939bae9c3700000000,
104'h5423794546d4196ca800000000,
104'h308d11401a16ec6d2d00000000,
104'h60c7849e8f1d7de33a00000000,
104'h30e3f082c73ea7f37d00000000,
104'hb8a435404872caf7e500000000,
104'h302fbd3b5f106ee92000000000,
104'h00b296bc65645bc1c816f27e2d,
104'h66c5d8da8b49c0cf9300000000,
104'h08a70b584eaec3205d00000001,
104'h2cf90988f26f8adfdf00000000,
104'hbc3b98257795a7ae2b00000000,
104'h2c07a6350fc364128600000000,
104'h669cf0ea39d25fc8a400000000,
104'h901a828935628929c5780ba0f0,
104'h940644390cb24d8a6400000000,
104'h30409af3818a989c1500000000,
104'h5457c759afc0fad08100000000,
104'h3013809d27c00eaa8000000000,
104'h943402576819f5353300000000,
104'h08708573e152814fa500000000,
104'h30efdc00df3e6a177c00000000,
104'h0872a823e57a9c45f500000001,
104'h346165e1c20a828f1500000000,
104'h94994016320ddd091b00000000,
104'h28596845b2267f7d4c00000000,
104'h00c7697a8e840ed4084b784e96,
104'h3053ae37a70f95791f00000000,
104'h2888313c10ca86a69500000000,
104'h54aa1182549488e02900000000,
104'hb8c3810687211f3d4200000000,
104'h945646b7ac6209d1c400000000,
104'h94cfcb469ffcf50ef900000000,
104'h300e691d1cfad024f500000000,
104'hbc8c772618ace25a5900000000,
104'h284846c1903777776e00000000,
104'h34f10c92e23bbb1d77ffffffff,
104'h086f6c71de2a1b275400000000,
104'hb83d20397acc490e9800000000,
104'h0459f1b7b301b24d0300000000,
104'h28b4ff82696b07b1d600000000,
104'h30c804e090492bc99200000000,
104'h94971c9c2e11a03b2300000000,
104'hbc7a36f7f49e4a323c00000000,
104'h28b63a746c5825adb000000000,
104'h902a87cb55bc3fe87896b8232d,
104'h08e458b4c81010bf2000000001,
104'hbc7431e3e8760b07ec00000000,
104'h661a5fcb34c4fbee8900000000,
104'h3476368fecfc9166f900000000,
104'h2c088ce111df1f78be00000000,
104'h90bca9da798c7ca81830d57261,
104'h947b9de3f7e38d58c700000000,
104'h9cbcbe90795fd627bf1c960039,
104'h60c2bd7e850e2d4b1c00000000,
104'h2cef923cdf7f62fbfe00000000,
104'hbc022f1f044178c98200000000,
104'h9c57b92bafcfc0029f4780028f,
104'h301ebaf13d07f7130f00000000,
104'h60fd8a68fb763dddec00000000,
104'h9cadd9dc5b2379214621590042,
104'hbcae2bc05c717ce1e200000000,
104'h2c16a1952de615b2cc00000000,
104'h2c095dc11201c92d0300000000,
104'h00cf707e9e50e541a12055c03f,
104'h30aa07b2543d369b7a00000000,
104'h946459cbc8b47e086800000000,
104'h08f583a2ebeb7ccad600000000,
104'h28b25164644f30079e00000000,
104'h90ddaa5ebb8593160b583948b0,
104'h668317f4062500f54a00000000,
104'h94a19f7043f50c98ea00000000,
104'h5475e6ebeb0d68531a00000000,
104'h00595d27b26f342fdec8915790,
104'h54e0dc72c1b2cb586500000000,
104'hbcd8008ab087e8760f00000000,
104'h301727772effb906ff00000000,
104'h0030d569615837c9b0890d3311,
104'h603ff3a37f35e6156b00000000,
104'h2ceb224ed654bc43a900000000,
104'h54aa156254aae9005500000000,
104'hbcb0b486612fb7bf5f00000000,
104'h9c4875e590e6b606cd40340480,
104'h30032c1d06e2efdcc500000000,
104'h60c33f14869fdb223f00000000,
104'h604407df88bd49f67a00000000,
104'h9c49c79b93d17c10a241441082,
104'h081b7157361027272000000000,
104'h34113ee922e70e4ace00000000,
104'h0809c8d313d8804ab100000000,
104'h602c192558b9d5107300000000,
104'h9caff15a5f7fc1ffff2fc15a5f,
104'h00263b3f4cdc1d5ab802589a04,
104'hb81a5cc1349068a02000000000,
104'h3091e6e0236e39e7dc00000000,
104'h941ad78b35fa5c46f400000000,
104'h60716679e2793f33f200000000,
104'h2c7d1509fa430cd38600000000,
104'h00297931528b7f7616b4f8a768,
104'h28a1fb4643bd4dde7a00000000,
104'h66687ef5d012c6af2500000000,
104'h08cdaf0e9ba4f2c64900000000,
104'h002e64735cb0569a60debb0dbc,
104'h28345fed68ba2aa47400000000,
104'h00e14f14c282a2b40563f1c8c7,
104'h3491d42c23b89c5671ffffffff,
104'h2c1b09073620cc374100000000,
104'h08d7b4dcafc642788c00000000,
104'h309b2d3636c3de208700000000,
104'h9c3e99c77db607666c3601466c,
104'h088a134e14d9c92ab300000001,
104'h08c5d5788bba213c7400000000,
104'h08f87bbcf0fe1fd2fc00000001,
104'h54ee013cdce22dd6c400000000,
104'h0847fbab8f1492552900000000,
104'h343a491f74810ed00200000000,
104'h94e82904d0012aad0200000000,
104'h60c477ec88568585ad00000000,
104'h00948678293a489774cecf0f9d,
104'h2cefc330df188f133100000000,
104'h94ff2f70fe305d8d6000000000,
104'h340657390cb880527100000000,
104'hb8944418284768cf8e00000000,
104'h664da30f9b7fe1e3ff00000000,
104'h90c2155e84de3354bc1c260a38,
104'h30dd647ebae10c1ec200000000,
104'hbcf210ece49f4bdc3e00000000,
104'hbc4574178a9783222f00000000,
104'h541e6d313c17c2e32f00000000,
104'hbcce51209c7412cbe800000000,
104'h30b09554614fa6a39f00000000,
104'h90e06da8c0f0aab2e110c71a21,
104'h3014554528e03f18c000000000,
104'h90de3a7cbc67fa35cfb9c04973,
104'h342bc5af57c40a008800000000,
104'h307cf327f98ccc701900000000,
104'h348ff7fc1fdc76d6b8ffffffff,
104'h306829f5d07d243ffa00000000,
104'h9c4a625d94e962d4d248625490,
104'h9cbc13f0788d183c1a8c103018,
104'h60730bb7e66e54f9dc00000000,
104'h9ca294e645a56ec64aa004c640,
104'h90df77bcbec17a00821e0dbc3c,
104'hbc1f0b633ed1f9f8a300000000,
104'h60ce52d49c4060658000000000,
104'h00d4dcb2a95bb3afb730906260,
104'h9c3bde2f77667463cc22542344,
104'h2c54c0e3a98a99841500000000,
104'h904b1bb596413bf7820a204214,
104'h543ccebd79eb48d4d600000000,
104'h00efba14df7e52dbfc6e0cf0db,
104'h2c3747cd6eb45abe6800000000,
104'h2cc4c0b8890f268f1e00000000,
104'h54a4245e48a7801a4f00000000,
104'h60bbfbce771e724d3c00000000,
104'hbc795f81f28a5d861400000000,
104'hbc12284124d37b0ea600000000,
104'h60a602fc4c13275f2600000000,
104'h2cb3dfba671f0b933e00000000,
104'hbc03f36107e4fdbec900000000,
104'h90ff44a8fe8e30541c7174fce2,
104'h04a47bf648f80882f000000000,
104'h048e6e381cdeb390bd00000000,
104'h60039acd078953461200000000,
104'h28769457edd15942a200000000,
104'h546e0cabdc6e6965dc00000000,
104'h2827fbab4f75db27eb00000000,
104'hbca619204c68b1fdd100000000,
104'h94daa1a4b5eca4b6d900000000,
104'h30931e7a26d48be6a900000000,
104'h2833a871675a4f33b400000000,
104'h0887ddc20fd029c0a000000001,
104'h288f82f81f88dd921100000000,
104'h046b86c5d7b62de66c00000000,
104'h001ce0e93972b897e58f99811e,
104'h08d1840ea38806741000000000,
104'h00b45aae68b36ab66667c564ce,
104'hbccc06ea98a409464800000000,
104'h9418dd73319a1c303400000000,
104'hbc0553650ae34ff8c600000000,
104'h600cd7271959cf01b300000000,
104'h546bcc4bd7fb53e4f600000000,
104'h66682273d0935ae02600000000,
104'h607cbf27f9bf4a2a7e00000000,
104'h341ab2c3353529516a00000000,
104'h00f9f046f39d3fa23a972fe92d,
104'h9cc80042906cb189d948000090,
104'h0495e6b42b72f4ebe500000000,
104'h9c6733e1ce25b4894b2530814a,
104'h00e2f83cc5967a5e2c79729af1,
104'h5414134728533909a600000000,
104'hb891156c22ae8c1a5d00000000,
104'h90fcace2f9fe4786fc02eb6405,
104'h94c6558e8cb6adfa6d00000000,
104'h6017c3df2fd6663eac00000000,
104'h901e42af3c4b079b96554534aa,
104'h9c0ffc271fbfd52c7f0fd4241f,
104'h309be59a371800553000000000,
104'h548fc6681f9b8a0c3700000000,
104'h049a91dc35099b491300000000,
104'h94da0c0eb444ec598900000000,
104'h608971c01296934e2d00000000,
104'h905b9b45b781515002daca15b5,
104'h00fdd254fb4337058641095a81,
104'hbca152f8425d37edba00000000,
104'h34682f65d03804c77000000000,
104'h00df0ed4be3344eb661253c024,
104'h5477ff79ef8806b01000000000,
104'h34f35346e658fec9b1ffffffff,
104'hbcfa3fe0f482ee9e0500000000,
104'h0093b978272d49bf5ac1033781,
104'h00bec0a87d2ef22d5dedb2d5da,
104'h900e1b571c04a3c9090ab89e15,
104'h60d03098a0c666b48c00000000,
104'h2cca7f8e942f20a75e00000000,
104'h940ae94315d51d56aa00000000,
104'hb879c58bf31425d32800000000,
104'h2cde7aecbc517eeba200000000,
104'h2c9d11763a1fe6873f00000000,
104'h34c5f8a68bcd680e9affffffff,
104'h54d1f840a3fe9fc2fd00000000,
104'h08c3043a869ac51e3500000000,
104'h540f6b951e61943fc300000000,
104'h2ce79a36cf7fee37ff00000000,
104'h34bf65da7e49c87993ffffffff,
104'hbcba9de47557c333af00000000,
104'h9c615643c2947eac2800560000,
104'h0403255106b987ac7300000000,
104'hbc214cb7424572d78a00000000,
104'h664685498d847f040800000000,
104'hb88fe5e41fcad6b29500000000,
104'hb8051d570aeb4852d600000000,
104'hb866f737cd370dbb6e00000000,
104'h0081e3c8035afa77b5dcde3fb8,
104'h5406fadb0d2c292f5800000000,
104'h30a0b1a8415a0009b400000000,
104'hb8193bb932f52406ea00000000,
104'h08274ec34e3ab3677500000001,
104'hb882c1820508df011100000000,
104'h2c6d3da5da3dbaad7b00000000,
104'h9493fc9e27f2dc98e500000000,
104'h284647998c8023b60000000000,
104'h2821323d425dbd0bbb00000000,
104'h08b3c8aa67d1401ea200000001,
104'h30efa848dfbb7a527600000000,
104'hb8a8bba8514c41459800000000,
104'h90a3916a47c7642c8e64f546c9,
104'h66ec861cd9519441a300000000,
104'h341ab91335dddc14bb00000000,
104'h54e88452d13bfdf37700000000,
104'h30dfef6cbfe5d144cb00000000,
104'hb8ec5558d8ed76f2da00000000,
104'h2c2335634647fcbd8f00000000,
104'h5434e6fb690fc79f1f00000000,
104'h0062a8a1c52fdd355f9285d724,
104'h08c241c084a4e4124900000000,
104'h30b02f926012732b2400000000,
104'h34c814fa9043082b86ffffffff,
104'h043fe5677f36bcdb6d00000000,
104'h904502b58a189381315d9134bb,
104'h04ab460856bbf2407700000000,
104'h9c0cabb71993a5742700a13401,
104'h28151a212a598117b300000000,
104'h28507b93a049791f9200000000,
104'h2c1a232134d4c8dca900000000,
104'h2c73348fe679815ff300000000,
104'hbc3a872f75e896ccd100000000,
104'h28b33bba664844cd9000000000,
104'h0827fd3b4f1a61e13400000000,
104'h08f7a4e0ef8df9c61b00000000,
104'h2824b8ef49b946d67200000000,
104'h2ccbfe8e97d4e268a900000000,
104'h945f16b9be02c42b0500000000,
104'h3456de0fade3688ec600000000,
104'h08f607c2ec2936195200000001,
104'h34d72b6caeedf9d2dbffffffff,
104'h08123df924b8129c7000000000,
104'h04f42d76e84ca3959900000000,
104'h2c4018098091e5722300000000,
104'h9cec55b6d8506eeda04044a480,
104'h94f64d5cec840c160800000000,
104'h086ecc7bdd947cba2800000000,
104'h2cf55a20ea2c31c35800000000,
104'h60abbccc57e6e196cd00000000,
104'h04ebab42d7ab8b745700000000,
104'h94e76078cea541de4a00000000,
104'h008a8a6c1563d3ebc7ee5e57dc,
104'h309bcc0c37292daf5200000000,
104'h30f7ca0cefba079c7400000000,
104'h08f57ad2eaa03ce24000000000,
104'h2c48314d909ae0c83500000000,
104'h54369ad76d6beb15d700000000,
104'h906ea819dd3d136b7a53bb72a7,
104'h304d18e79ae533a4ca00000000,
104'h94cc231e985d493dba00000000,
104'h28a76c8c4e1fedab3f00000000,
104'h604c4fc998efddbedf00000000,
104'h041424172809e8071300000000,
104'h94bb004276045a290800000000,
104'h6638308d7001c5510300000000,
104'h34be577a7c56b17badffffffff,
104'h30e7f1c0cfc197e68300000000,
104'h08a1b51a43ca3c6c9400000001,
104'hbc6f0239de393de57200000000,
104'h66dd6190baca757c9400000000,
104'h3092c34425b47d246800000000,
104'hbc06fa070d4d74e79a00000000,
104'h00dba8f0b768df47d144883888,
104'h28969c682df42ca6e800000000,
104'h54714607e2474da58e00000000,
104'h30acd364598464780800000000,
104'hbc9518122aad6d585a00000000,
104'h08c542648ab875d67000000000,
104'hbc8813601052bb41a500000000,
104'h660211970420c8014100000000,
104'h3066eeffcd8d67fa1a00000000,
104'h2c7c19e3f8930bee2600000000,
104'h084930b792caf3de9500000000,
104'h60c3d0fa87633861c600000000,
104'h94aef9165dd88b0ab100000000,
104'h047ef545fd6245cfc400000000,
104'h28098f6913572159ae00000000,
104'h94cef9f09d5eaa77bd00000000,
104'h08eaadb8d5774e69ee00000001,
104'h2cec32ead8a296544500000000,
104'h28268cd54dd8e994b100000000,
104'h3021c0db43abef225700000000,
104'h00f4b046e92a65f7541f163e3d,
104'h66163d312c1a0c613400000000,
104'h08db725cb6e3ee6cc700000001,
104'h9c0d26191a8d33461a0d22001a,
104'h60f25020e43a41957400000000,
104'h008d0a7c1af3d2d4e780dd5101,
104'hb8c6f55e8d254dc74a00000000,
104'h2c9676082c817fc20200000000,
104'h04f108a4e2168d212d00000000,
104'hb8579d29af4bb08f9700000000,
104'h5420b73d41bb217c7600000000,
104'h6008c90b114839759000000000,
104'h2834013368e5b07acb00000000,
104'h545d839bbb2988715300000000,
104'hb89ec5543d7bff75f700000000,
104'h66b683806d54a13fa900000000,
104'h90318d2d63044f850835c2a86b,
104'h2800582f00ecd958d900000000,
104'h9c0b1909162e79895c0a190914,
104'h90ead5cad5b153fe625b8634b7,
104'h6040abf18174ca1de900000000,
104'h9ce54144ca283e295020000040,
104'hb88917b612b09d9e6100000000,
104'h900b3c471653ca95a758f6d2b1,
104'hbcf688e0ed3ebc257d00000000,
104'h90ee713edcecedc0d9029cfe05,
104'h908b12be160f75911e84672f08,
104'h9ce8ff56d1dfd9e4bfc8d94491,
104'h9433fb5d67be7d7c7c00000000,
104'h0464a67bc9863afc0c00000000,
104'h6677c785ef8e87441d00000000,
104'h2c42b35985db32c8b600000000,
104'h04e306c2c6e4a202c900000000,
104'h2850ab5ba1a514c24a00000000,
104'hb8ffdf62ff9f54943e00000000,
104'h0875b8adeb50e225a100000000,
104'h28645a73c8657997ca00000000,
104'h9004d63d09fb85eef7ff53d3fe,
104'h04236fbd46c8db649100000000,
104'hbc5fbbb5bfe4d0d8c900000000,
104'h94acd1ce59d8901ab100000000,
104'hb8d68982ad4835619000000000,
104'h90e779f2ce7f1595fe986c6730,
104'h087034d1e05743c3ae00000000,
104'h0012f43525c82d6e90db21a3b5,
104'h2c07b38b0fd1e5faa300000000,
104'h30bb6b6276ea7902d400000000,
104'h04e9e85ed3785bc5f000000000,
104'h66cc750698b0d5706100000000,
104'h28e04eb6c052f69ba500000000,
104'h548e9d6e1d9f77903e00000000,
104'h945466bfa88b95bc1700000000,
104'h041bb3a537f0c800e100000000,
104'h90f7e164ef54e223a9a3034746,
104'hb895d5742b45ff1d8b00000000,
104'h041d8c533b1b4a8b3600000000,
104'h342d3b6d5aa781004f00000000,
104'h60aefdf65dfbbf70f700000000,
104'h30c0c4d68130f9896100000000,
104'h906b017bd63c2f1178572e6aae,
104'h66a543be4a8538500a00000000,
104'h28d8c2cab141c1678300000000,
104'hbcdf88f2bfe5ccb2cb00000000,
104'h341bba953740d42f8100000000,
104'h04dd2ffcba8a61ce1400000000,
104'h28945a4228a2b6e44500000000,
104'h08782b2bf093da7c2700000000,
104'h08f97802f2dd26c2ba00000000,
104'h66d10f86a2b72d5a6e00000000,
104'h30567abdac378ac76f00000000,
104'h664c20dd987c00c5f800000000,
104'h301a462334b9efae7300000000,
104'h2cbd1db87aab06d65600000000,
104'h0022e69b4541c3f38364aa8ec8,
104'h308dcb681b48196d9000000000,
104'h0871fd55e37853d1f000000001,
104'h346b41f9d63416236800000000,
104'h9cf5ec3aeb2705454e2504004a,
104'h9cc5f8328b527a53a440781280,
104'hbc93c1fa272554094a00000000,
104'h34308fa361cebf1c9d00000000,
104'h605de5ffbbdc8d9cb900000000,
104'hb8696095d2dd7558ba00000000,
104'h9ca38474471d4d3b3a01043002,
104'h349ac616351521a52affffffff,
104'h0044ba4789c2b7dc850772240e,
104'h941e29f33c3ad85d7500000000,
104'h2c778121ef5f7841be00000000,
104'h28cdd0b69b1e999d3d00000000,
104'h2ce95b6ed2f07ae2e000000000,
104'h9cb165ac62e36d40c6a1650042,
104'h04e9c05ed35169ffa200000000,
104'h549146e222cf3ee49e00000000,
104'h660947dd12eee990dd00000000,
104'h04bc9120797e79e3fc00000000,
104'h04599691b3f29354e500000000,
104'h600debf71b17655b2e00000000,
104'h603a09eb74e4b2c4c900000000,
104'hb8fb15b0f6d94024b200000000,
104'h285d2417ba7fc121ff00000000,
104'h283b2f5976231cdf4600000000,
104'h9c72b7ffe531a1616330a16161,
104'h544fc8bb9fce7de49c00000000,
104'h30a2d54e45869c440d00000000,
104'h28fcac64f979b153f300000000,
104'h00c574748a7a1c45f43f90ba7e,
104'h947a6ba1f41ded053b00000000,
104'h0802e2990569299fd200000001,
104'h04efaa7adf0d2a971a00000000,
104'h9048edad9122a64f456a4be2d4,
104'h907d2bc1fa33c363674ee8a29d,
104'h30c0d05881514a0fa200000000,
104'h30e89cfcd139cc897300000000,
104'h9c31de09633b5e5f76315e0962,
104'h94b2227c64e032e0c000000000,
104'hbcfceee8f9943a762800000000,
104'h6620a34b41b597086b00000000,
104'hb81c8be739db7f56b600000000,
104'h9490d53221fee95cfd00000000,
104'h9455daadab8613b60c00000000,
104'h601308c3266fc5f9df00000000,
104'h088649a80cece014d900000001,
104'hb823b545470e90b91d00000000,
104'h9cb9fc0473bd4aac7ab9480472,
104'h2c0ac4c515605139c000000000,
104'h2876f5aded67737bce00000000,
104'h082da0115bb84ed27000000000,
104'h3069074fd2c6303a8c00000000,
104'h305ffab3bf476ca78e00000000,
104'hb85a7a55b4fcc866f900000000,
104'h28ff5ef6fe47458d8e00000000,
104'h34257ceb4a46713f8c00000000,
104'h046579ebca5d0823ba00000000,
104'h2c0a4dff143389bb6700000000,
104'h60fd275afa1012c52000000000,
104'h2896293a2c9096982100000000,
104'hbc063dcf0cf04f8ee000000000,
104'h2c06f30d0df2fe56e500000000,
104'h66d41a96a8c8505c9000000000,
104'h60d7a49eafa7852c4f00000000,
104'h5412edbf25f72acaee00000000,
104'hbce177dcc27e8917fd00000000,
104'hb85fc60fbfce14329c00000000,
104'h303dd3757bb1fdd46300000000,
104'h543f5d197e8dbdb41b00000000,
104'h90d4f6d0a9e128e0c235de306b,
104'h543fa3237f5f7029be00000000,
104'h9445661d8ade1d74bc00000000,
104'h00d00b3ca065e82dcb35f36a6b,
104'h9090164620c8f8909158eed6b1,
104'h541c973139c1f21c8300000000,
104'hb8b558fa6ab4dcec6900000000,
104'h28f7a38cef26c6154d00000000,
104'h302e88a15dd2af06a500000000,
104'h349e739a3c5a23f1b4ffffffff,
104'h28f07468e0dd911abb00000000,
104'h30e47d66c8bc2f4a7800000000,
104'h90628c3dc5451f258a2793184f,
104'h601175bf22b30b826600000000,
104'hb876cccbed516ae1a200000000,
104'h547e1c2dfc9637b02c00000000,
104'h30ce6b7c9c3cb7c97900000000,
104'h00bbc6fe7775aab5eb3171b462,
104'h309742802efef71cfd00000000,
104'h54d2af3ea5d8af26b100000000,
104'h908dfcbe1b4703d58ecaff6b95,
104'h66e2fcb8c5507f65a000000000,
104'h305101e9a2dd9eaebb00000000,
104'h283491fb697aa18bf500000000,
104'hbcf02264e06e2a27dc00000000,
104'h9c81984e03cf03749e81004402,
104'h90650363ca712679e214251a28,
104'h0807cbc10f55d6bdab00000001,
104'hb8604acfc0b46da06800000000,
104'h54ac871e59212cc34200000000,
104'h30978b502fbd2f5a7a00000000,
104'h083f8ff37f26529f4c00000000,
104'hbc7ff059ffffad22ff00000000,
104'hb8a8a28851d2ed30a500000000,
104'h9021aa1343a8b63251891c2112,
104'h088bbdee1779d511f300000001,
104'h28701969e074e38be900000000,
104'h04b02ff06073b29de700000000,
104'h9c52bc07a5d193e2a3509002a1,
104'h083661176c8f59f01e00000000,
104'h304ad8599543a7b98700000000,
104'h306860b1d02de6e95b00000000,
104'h2861e98dc3cffd489f00000000,
104'h54b130ca6226991f4d00000000,
104'hb8cccb8e99e1ac8ec300000000,
104'h2c06d22d0d4e6ff39c00000000,
104'h286fa707dfea0344d400000000,
104'hbcd31068a63f867d7f00000000,
104'h942e9d675db640ea6c00000000,
104'hbc270dc54ebc2f9c7800000000,
104'hbcb734d46e3712bb6e00000000,
104'h00c58f508bc9d1ea938f613b1e,
104'h002e84415d35cfaf6b6453f0c8,
104'h945008d7a05f83c5bf00000000,
104'hb8f01f54e03374856600000000,
104'h60a268e4444467478800000000,
104'hbc49c27f936d5fb9da00000000,
104'hb829a4c55379c64df300000000,
104'h08dfbee8bfc3cd868700000000,
104'h54c10482824cee719900000000,
104'h3026267f4cfe13eafc00000000,
104'h34622eedc4eccd12d900000000,
104'h661ab7ef35a89ea05100000000,
104'h2cb3f58c671f4b4b3e00000000,
104'h2c2b8aa35788ab241100000000,
104'h9443e0b1877269f9e400000000,
104'hbcf67ac6ec61c4b1c300000000,
104'h9cf67b62ec051db50a04192008,
104'h284d55499a8900421200000000,
104'hb8fa5f6ef4c3eadc8700000000,
104'h28aac3d25581f8980300000000,
104'h344a016394b5418c6a00000000,
104'h2803f8d307a18a2a4300000000,
104'h30883c8810b199a06300000000,
104'h60a31b7246724f37e400000000,
104'h28c39eec87a34eb24600000000,
104'h9076739fec56dbb9ad20a82641,
104'h9c6c755dd82a3c235428340150,
104'h5400560500a5b96a4b00000000,
104'h60899762133f19097e00000000,
104'h04d3d00ea73b23cd7600000000,
104'h28f7f34cef3294456500000000,
104'h9c4a13e9943c84177908000110,
104'h9c40da238124306f4800102300,
104'hb8dca480b989ad481300000000,
104'h34530bb7a6ccdfe49900000000,
104'h66504181a017d81b2f00000000,
104'hbc2a828f553960c37200000000,
104'h049c935639325f0b6400000000,
104'hbc32fffb65d058e2a000000000,
104'h603c972d795d3a55ba00000000,
104'h2cf15806e2c031e48000000000,
104'h9c53caefa7553bf5aa510ae5a2,
104'h043f7d7d7eb0b5226100000000,
104'h04d4194aa86a0ba7d400000000,
104'h90274de94e5467b7a8732a5ee6,
104'h089085aa212de2e55b00000001,
104'h34281d975035a67f6b00000000,
104'h04e8983cd13708ef6e00000000,
104'h34730395e6db8218b700000000,
104'hbc7889e9f16f0ebdde00000000,
104'h6069e5add3225add4400000000,
104'h04fa3060f42bcb0f5700000000,
104'h046d446dda643ce9c800000000,
104'h3442aa0b850e165d1c00000000,
104'h00c4c71e89ccfc169991c33522,
104'h9008ca17116246e5c46a8cf2d5,
104'h542e87cf5df61006ec00000000,
104'h04e04470c07e6ca3fc00000000,
104'h9c611f4bc2a630124c20100240,
104'h9c9599c02b5a4d51b410094020,
104'h348c711c1850af55a1ffffffff,
104'h2cd6c376ad5d206fba00000000,
104'hbca537924ab098aa6100000000,
104'h04d49fbea91d0b353a00000000,
104'hb8074fb70e9b8ab23700000000,
104'h2c491d83928c5ca21800000000,
104'h28bac55475e853c4d000000000,
104'h600e286f1cd08970a100000000,
104'h00679efbcf054dff0a6cecfad9,
104'h283154ef62bee81c7d00000000,
104'h04c469f2889a7b3a3400000000,
104'h60304c3160bb2ce27600000000,
104'h600b864917536119a600000000,
104'h30c9f8209373a5bfe700000000,
104'h90c332ca86aca4f2596f9638df,
104'h00906f6620b7366c6e47a5d28e,
104'hbce45902c86167e3c200000000,
104'h6627a1754f611467c200000000,
104'h602c193f58d462c6a800000000,
104'h04dcc270b91642ed2c00000000,
104'h662416874890c23a2100000000,
104'h5402774b0450cef7a100000000,
104'h602d82ad5bbec29c7d00000000,
104'h043dc1ad7bf4cb42e900000000,
104'h309aea3635280c035000000000,
104'h54afac045f6b0c4fd600000000,
104'h08a4c0744927ce4f4f00000001,
104'h04a7b57c4ffda452fb00000000,
104'h90c4ab7289a29d1a45663668cc,
104'h664afe0195f21f4ae400000000,
104'h28c38ffa87e20bc2c400000000,
104'h005c323fb89d7ef63af9b135f2,
104'h94865d980cf00960e000000000,
104'h901037a1206df6d1db7dc170fb,
104'h30659a99cbcdfcd29b00000000,
104'h089b985237a668124c00000001,
104'h669bb00837a3a0b44700000000,
104'h08e4af42c9479dbd8f00000001,
104'h2c15f5b32bc19f628300000000,
104'h0486941a0d634887c600000000,
104'hb8b47e246813eef92700000000,
104'h9010c74921d4baeea9c47da788,
104'h54c4a2a8895fed53bf00000000,
104'hb82f9df75f1b65313600000000,
104'h9c424f4b846a3c0dd4420c0984,
104'h08296e1152d31148a600000000,
104'h302c0ed958e05c80c000000000,
104'h28dc7a44b805def30b00000000,
104'h94f5d6dceba20bce4400000000,
104'h34299dfd5353ffa9a700000000,
104'h30e693a4cdc65ece8c00000000,
104'h0077b965efad32aa5a24ec1049,
104'h90ec743ad8789e1ff194ea2529,
104'hb8bbdd6a771800f13000000000,
104'h3433f66b6788e21a1100000000,
104'h083237b964c2b9388500000000,
104'h908db2c21b4c6edf98c1dc1d83,
104'h28b3bebc675a2bffb400000000,
104'h306ee88ddd29d0475300000000,
104'h28549da1a962277fc400000000,
104'h2818c9d531ecb5eed900000000,
104'h60b760506e0bb3b51700000000,
104'h0432876965bd8f307b00000000,
104'h0840df7b81c50e5c8a00000000,
104'h94e21cd2c458e72db100000000,
104'h6618ec89317f66f3fe00000000,
104'h2c2fdc615fe280bac500000000,
104'h30a3bda847665ab1cc00000000,
104'hb840bb1d81703279e000000000,
104'h66e019c2c08530940a00000000,
104'h30b35cd2662882c35100000000,
104'h30d64488ac95d55c2b00000000,
104'h2c2be00f579103b42200000000,
104'h2803aa6107f59780eb00000000,
104'h00da6a1eb4686f2bd042d94a84,
104'hbc6f4c7bde7ba33ff700000000,
104'h9488730e102882c15100000000,
104'h94d2ecc0a5ad3e925a00000000,
104'h0078d1a9f10b9bd117846d7b08,
104'h9404f9e1098bc5361700000000,
104'h662687794d32137b6400000000,
104'h608f3b441ef864aaf000000000,
104'hb8ae4cca5c435a978600000000,
104'h901e3d1b3c699829d377a532ef,
104'hbc6edcaddda6d5c24d00000000,
104'hb8357c4d6a6e64abdc00000000,
104'h302c00e95830795b6000000000,
104'h28545287a83b54ef7600000000,
104'h00c05e0c80dd257aba9d83873a,
104'hb877a235ef3d35717a00000000,
104'h3429ff6353fac1fef500000000,
104'h60a44284486d906ddb00000000,
104'h9c7da2f9fbd81a82b0580280b0,
104'h66e62b62cce4e9dec900000000,
104'h9c0cc59719d87a60b008400010,
104'h00f06176e0e6bb82cdd71cf9ad,
104'h00ca6ecc948708b80e517784a2,
104'h2c49a231936330d3c600000000,
104'h30babce67505e4630b00000000,
104'h94b1cfbc63aaa30e5500000000,
104'h66f930eef2f4fffce900000000,
104'h542c1d0558ced52e9d00000000,
104'h54a1bab043acbde25900000000,
104'hb8d9f9b4b3edeff2db00000000,
104'hbca884ba51684c31d000000000,
104'h6092be3a25633dd3c600000000,
104'h666c8057d9bbc0c27700000000,
104'hbce417bec899a70c3300000000,
104'h6690b1902171f535e300000000,
104'h66e73432cefbed9cf700000000,
104'h2c683b37d0ae22e05c00000000,
104'h9c16ae3f2d3ea93d7d16a83d2d,
104'h00012ad302ed3ee6daee69b9dc,
104'h0011394f2200036d00113cbc22,
104'h549a04b23443161f8600000000,
104'hbcf50d8eea793365f200000000,
104'h080e0fe11cef2926de00000000,
104'h66c013ec80bdba247b00000000,
104'h088462280825485b4a00000001,
104'h60e0d212c1c45e648800000000,
104'h306dac19dba5efd64b00000000,
104'h9ce4166ec835e8a36b24002248,
104'h289cc4fa398263760400000000,
104'h30eb642ad6bd9f1a7b00000000,
104'h0005f6db0b288ad7512e81b25c,
104'h00581f33b05781c9afafa0fd5f,
104'h9c710a87e2928d502510080020,
104'h08d77834aed84668b000000001,
104'h342a138954362e056c00000000,
104'h9cbb189a76ab147456ab101056,
104'h547cfc2df90fe7cb1f00000000,
104'h664a8e919581012c0200000000,
104'h6087d1800fe5c940cb00000000,
104'h04797905f26e4b89dc00000000,
104'hb8afcf505f9e10c23c00000000,
104'h302e73a15cb158466200000000,
104'h00c52c248a45886d8b0ab49215,
104'h3406c2d30d1f6de53e00000000,
104'h66a1a54c4321a21b4300000000,
104'h2842bfc585f3309ae600000000,
104'h08cdcad49bea5368d400000001,
104'h084704638e78de65f100000001,
104'h60790b85f207b1b10f00000000,
104'h34de575abcd44b02a8ffffffff,
104'h08d080eea16f4e13de00000001,
104'h6628581750dc9beeb900000000,
104'hbc807b58007d5167fa00000000,
104'h94e0eac2c1c9c4629300000000,
104'h34eccdd2d9e5584acaffffffff,
104'hb86c644dd82fc15f5f00000000,
104'h306bda27d7970f1a2e00000000,
104'hb8d47660a883959a0700000000,
104'h94905ce220328df36500000000,
104'hbca1db66432605954c00000000,
104'h664df9519b6874afd000000000,
104'h343ec28f7db013886000000000,
104'h9484857c0961c6e9c300000000,
104'h284dfbc39bfd3b72fa00000000,
104'h603e16357c0b88011700000000,
104'h6622e3b1452f6f0f5e00000000,
104'h2cabcb0257e2170ec400000000,
104'h08460fc38ca8d1d65100000000,
104'h04ad5a345a984af23000000000,
104'h28b2ba2665b7350a6e00000000,
104'h086f5cd5deb64e446c00000000,
104'h9038edc5716d53a3da55be66ab,
104'h006c5aafd80c3b6318789612f0,
104'h6630724f60e5ce5ccb00000000,
104'h04dc9650b99478682800000000,
104'h5468782bd0ebe7b4d700000000,
104'h30609905c121d3334300000000,
104'h9000048900c5ffe68bc5fb6f8b,
104'h00727ed7e4f55d5aea67dc32ce,
104'h2c931d54269dd0ee3b00000000,
104'h54ea0294d41808413000000000,
104'h04e8b536d1c26a888400000000,
104'h909f49c83e1400fd288b493516,
104'hbc0d579f1abfee307f00000000,
104'h90f870bef069cc6fd391bcd123,
104'h9c8694b80d090b211200002000,
104'h60edd684dbdd232eba00000000,
104'h040b2d6f16ae3a585c00000000,
104'h60d128e6a2758d9beb00000000,
104'h2cebff6cd75eba91bd00000000,
104'hbce3306cc6cebfce9d00000000,
104'hb819b11f33af4c465e00000000,
104'h94845c660814b5a72900000000,
104'hb8731db3e662adb7c500000000,
104'h608c0ee018c78ebc8f00000000,
104'h90c88114912fd6dd5fe757c9ce,
104'h0812a8a325232a714600000001,
104'hbcbf63ec7e41f5738300000000,
104'h66ba553e74c683da8d00000000,
104'h9c8347ac066e28f9dc0200a804,
104'hbc4296fb85f6cddaed00000000,
104'h54ef127adedafea8b500000000,
104'h08f292e6e59a4f083400000000,
104'h049b3b463695ad7c2b00000000,
104'h2c261ccd4cc6fdc28d00000000,
104'h66fcb5baf9511233a200000000,
104'hbc09833b1380dc240100000000,
104'hbc809e44014a6b479400000000,
104'h08501b7ba004140b0800000000,
104'h3450a60fa10fd4f51f00000000,
104'h94718d99e3b6d30e6d00000000,
104'h902c3f0558a485384988ba3d11,
104'h90b9e062739ee6903d2706f24e,
104'h2c8287d4053ec7cf7d00000000,
104'h3438456370f717a8ee00000000,
104'h54b8f7e8719bba323700000000,
104'h6658a4e7b14047378000000000,
104'h9c4acb6d95a4c79e4900c30c01,
104'h28b3e9f867ea49d2d400000000,
104'h342d2f4f5ae2e510c500000000,
104'h00630e65c67083dbe1d39241a7,
104'h90a42d3848fb8d46f75fa07ebf,
104'h08e0e6b8c186456a0c00000000,
104'h34745799e8337cb96600000000,
104'h5446ae3f8daee65e5d00000000,
104'hb81d35993ab32da46600000000,
104'h906f5303de5da251bb32f15265,
104'h30886f24100914071200000000,
104'h604d81d39b7934a1f200000000,
104'h9059b8ebb32599994b7c2172f8,
104'h3480723800df3466beffffffff,
104'hb8cb805497ccd9da9900000000,
104'h00f37282e64330838636a3066c,
104'h00c4578e883a1e0574fe7593fc,
104'hb81433b928858b8c0b00000000,
104'h9491218622711917e200000000,
104'h08ebd5acd75e17e3bc00000001,
104'h946ffde7df78e3c9f100000000,
104'h5426b2e54df673a0ec00000000,
104'hbcd7f51caf7cb899f900000000,
104'h9cd6ecb0add024a0a0d024a0a0,
104'h66296453528e6fc21c00000000,
104'h667db71dfb1274832400000000,
104'h2c3329756686bb420d00000000,
104'h00a764f24e1c0ca138c3719386,
104'h9cb88f30713f22d57e38021070,
104'h662633bf4cf45214e800000000,
104'h66e3f8f0c721bff34300000000,
104'h60b7d7cc6ff881bcf100000000,
104'h90524ee3a4cab9dc9598f73f31,
104'h28a1c82a43e08c36c100000000,
104'h002329ef4637818b6f5aab7ab5,
104'h54904aa220f7b1daef00000000,
104'h2839bfc773bfcdbc7f00000000,
104'h90c43fc28824dec749e0e105c1,
104'h089a8ed035d456eaa800000001,
104'h945baed5b71ec6d53d00000000,
104'h3491ca3c233f53537effffffff,
104'h604111e582e7c1a4cf00000000,
104'hb80e85f71d62b2f1c500000000,
104'hb80d61c11a6d6691da00000000,
104'hbc5ea2a7bdb01b7e6000000000,
104'h94e8e1f2d1e7e8b2cf00000000,
104'h543779bd6e56a47dad00000000,
104'h2836acc96d5532e9aa00000000,
104'h90b749646ee25322c4551a46aa,
104'h6696ff4c2d2bc3d15700000000,
104'h90cb608896495671928236f904,
104'hbc8c454a182149c34200000000,
104'h04270ad54ea3031e4600000000,
104'h08cee5509da0fedc4100000000,
104'h00b73cb46e848faa093bcc5e77,
104'h041bcca9374dc4f99b00000000,
104'h543eff577dbf90507f00000000,
104'h0009bb5f13ac01b658b5bd156b,
104'h04889ca611fe330cfc00000000,
104'h9031504162cf3a709efe6a31fc,
104'h94578b4daf793b9bf200000000,
104'h04b3d4d867a770404e00000000,
104'h30071abb0ec3bf748700000000,
104'h34ecc974d94a3c0594ffffffff,
104'h3481df160368a1dbd1ffffffff,
104'h2cda311cb453aa59a700000000,
104'h94fddd50fbd5cfc4ab00000000,
104'h2c879da20f3ad79b7500000000,
104'h30a9771252d13bf0a200000000,
104'h3487fb8c0f364be16cffffffff,
104'h603516cb6a739adde700000000,
104'h344a1e2b940c170d1800000000,
104'h08e59ba2cb64dec1c900000001,
104'h94d40b88a8e9acb8d300000000,
104'h289b858637d67398ac00000000,
104'h2c310871621f80413f00000000,
104'h2cfae124f5773b25ee00000000,
104'h289e646e3c5c60bfb800000000,
104'h669ff3e63f5d48dfba00000000,
104'hbc4305cf86c495108900000000,
104'hb80ca7f919a15e004200000000,
104'h30fdb59efb00b7d30100000000,
104'h94bab8487528258b5000000000,
104'h08962ba82c2053614000000001,
104'h947e9c81fdd53034aa00000000,
104'h9c5cda7bb9ec3dd6d84c185298,
104'h3027350f4e23b07d4700000000,
104'h28057b5f0a04b5110900000000,
104'h3006371d0ce0f69ec100000000,
104'h54485a6190e73aaace00000000,
104'h54cd58969a84ac960900000000,
104'h5496624e2cb82ffe7000000000,
104'h60ec3c2ad862d221c500000000,
104'h28ebe8b2d76c322dd800000000,
104'h605b1d43b6b378b66600000000,
104'h9c8e39da1cad360c5a8c300818,
104'h667e3c0bfc2c3f995800000000,
104'h663fe4d17f97643c2e00000000,
104'h948e09701ca78fbe4f00000000,
104'h6637c7616f29b5195300000000,
104'h04b0131e601597e72b00000000,
104'h2ce6da18cd064cbd0c00000000,
104'h66acaf8259b3088c6600000000,
104'h9058bc43b1de9704bd862b470c,
104'h94ed69c6da418fed8300000000,
104'h54baffea75a7238c4e00000000,
104'h54302dd760be16027c00000000,
104'hbc5735dfae6f41afde00000000,
104'h601b346136d0b88aa100000000,
104'h900bb9a917785c8bf073e522e7,
104'h9c9daece3bf28700e590860021,
104'h340f3d971ee916f8d200000000,
104'h04c9334e9204fe9f0900000000,
104'h088b16b2163827977000000001,
104'h608fe8c81fd74662ae00000000,
104'h285848c9b02af4c15500000000,
104'h049372ee26d52b0aaa00000000,
104'h28eb5264d603f0930700000000,
104'h2cf09e26e1dbdb0eb700000000,
104'h283ab8d5753cb4e97900000000,
104'h66b3cba067f062ace000000000,
104'h9c2c542558e7df5ecf24540448,
104'hbc621d47c453e7e1a700000000,
104'h60d55b1eaa96ad4e2d00000000,
104'h94c361c68631a6656300000000,
104'h60992f4e325e57d9bc00000000,
104'h08d8c08ab1e2abb8c500000001,
104'h9cf2e900e5592fd5b2502900a0,
104'h9cac25c0588353160680010000,
104'h5475a343ebbf79e07e00000000,
104'h30646e53c8568179ad00000000,
104'h904f87df9f740a59e83b8d8677,
104'h9cca53ec9432a19d6502018c04,
104'hb85b9b63b7a0a1584100000000,
104'h002a18fb54f45ffee81e78fa3c,
104'h088e49181cbe06bc7c00000001,
104'h663df4ab7bb326da6600000000,
104'h6648af0f9123e6214700000000,
104'h008d3ee81a335a2d66c0991580,
104'hb8deaa0cbdfc6adef800000000,
104'h306c5c5dd8d253b0a400000000,
104'h905ba1a3b7379c176f6c3db4d8,
104'h9c896a7612e81ee0d0880a6010,
104'h6652141da4da78a0b400000000,
104'h60b1ab62635af4fdb500000000,
104'h3041e28583c5d31a8b00000000,
104'h603bb20b77e078fcc000000000,
104'h94e15ca6c2d0ede0a100000000,
104'h54424e1b8428b3a15100000000,
104'h94550d11aad3d70ea700000000,
104'h349c380038eecf60ddffffffff,
104'h2c22450d44fd8480fb00000000,
104'hbc3c7ce578ab947a5700000000,
104'h606868a7d091afd22300000000,
104'h9c67aab9cf65a4ebcb65a0a9cb,
104'h08acfaac59ea725ed400000001,
104'h30e9bc24d3db786ab600000000,
104'h664668a98c59a145b300000000,
104'h0438c4957103187b0600000000,
104'h903196e96345e95d8b747fb4e8,
104'h08305c35609b9c523700000000,
104'h28de2c76bc9fab443f00000000,
104'hbcd1cbf2a34c64f39800000000,
104'h663d9f1f7b8997581300000000,
104'h0034f979698e19121cc3128b85,
104'h6020ff6f41d109b4a200000000,
104'hbc9613342c596131b200000000,
104'h54b184b0639226342400000000,
104'h542bfc5157576389ae00000000,
104'h348fd8f01f23b47547ffffffff,
104'h943378b9661000172000000000,
104'h2ce624fccc26bbcf4d00000000,
104'h085b191bb651cc97a300000000,
104'h3478dc5ff155df63ab00000000,
104'hb87be6e1f7cfd0829f00000000,
104'h3482496204707a09e0ffffffff,
104'h2c4ad03795b1011a6200000000,
104'h54e4d916c95d7a5fba00000000,
104'hbc6ed40bdd8d7d561a00000000,
104'h340027470061fec1c300000000,
104'h9c27ee074f1589f52b0588050b,
104'hbc34ca7b6907b14b0f00000000,
104'h6072c299e55e4d73bc00000000,
104'h2ce2e002c50ee3d91d00000000,
104'h90550aebaa904c0820c546e38a,
104'h2c6f57ebde886c061000000000,
104'hb8bec0e87d73a3b3e700000000,
104'h609c00fa38f33f2ee600000000,
104'h2c2c0b41581608312c00000000,
104'hbc3e54c57cf9ce70f300000000,
104'h94f3e95ce7867efc0c00000000,
104'h3021038f422b22a55600000000,
104'h28ef9f68df62db51c500000000,
104'hbc9c406838cbb8689700000000,
104'h94e6e252cdb2fa2c6500000000,
104'h2c30cd1d619a1c183400000000,
104'h90ecc3c6d94dbe499ba17d8f42,
104'hb831c639632345d14600000000,
104'h9c995e2c32c3cc2287814c2002,
104'h66492f079202b56d0500000000,
104'h60cc40b4988c05f61800000000,
104'hbc633d93c62a4e875400000000,
104'h08639b49c7edc7c0db00000000,
104'h304c66ab980df47f1b00000000,
104'h00142a9728e4e33cc9f90dd3f1,
104'h940e29d91c4ee66d9d00000000,
104'h544de4099bfb5be4f600000000,
104'h9cd69d6aad42db318542992085,
104'h28d961ccb2d4e2f8a900000000,
104'h28f6ba6aed72dd63e500000000,
104'h949a0eca34e81370d000000000,
104'h004368a586ede760db31500661,
104'h30a112b442a16e0a4200000000,
104'h04e54aa6ca0b3f471600000000,
104'hbc7cfdf1f9ec1542d800000000,
104'h346349bbc6f892f0f100000000,
104'hb87235afe4dc4954b800000000,
104'hb873e1ede72fd3f95f00000000,
104'h90081fdb10f7a43cefffbbe7ff,
104'h28e12e0ac2b0d3be6100000000,
104'h34170f1d2e5715b7ae00000000,
104'h9c8bb39e179a9f5a358a931a15,
104'h5442eee5859e9f3e3d00000000,
104'h9057eef5af809bac01d77559ae,
104'h088eaf5e1d86d00e0d00000000,
104'hb8929f1a2597614c2e00000000,
104'h30747175e8740127e800000000,
104'h6617d1dd2f9558982a00000000,
104'h00ae72d25c57513fae05c4120a,
104'hbc48afc391e315acc600000000,
104'h349cb9e439d560d4aaffffffff,
104'hbc9c081c38777465ee00000000,
104'hbcf381d8e76ece25dd00000000,
104'hbc559cf7ab7b745bf600000000,
104'h2c1e669b3c26712b4c00000000,
104'h28b02f186091d4ee2300000000,
104'h348450d208e157a0c2ffffffff,
104'h08864a140c5e7139bc00000001,
104'h2c9821f2307c8107f900000000,
104'h0445d0318ba95c185200000000,
104'hbc622021c4545a97a800000000,
104'hbcba467c7439bc277300000000,
104'hb8ee224cdcb9fb4a7300000000,
104'h90f9e0c2f34467c188bd87037b,
104'h9cca7c2094921fe024821c2004,
104'h34814d90020a410314ffffffff,
104'h9083aa0a0719e6d5339a4cdf34,
104'h084a4231940251c90400000000,
104'h34c8bd34918d4c621affffffff,
104'h6068c6afd1aba7ac5700000000,
104'h30a4878a492b66875600000000,
104'h047b41d9f6e2f00ec500000000,
104'h60f787baefd460fca800000000,
104'h90f94538f257d407afae913f5d,
104'h541e952f3d3d39417a00000000,
104'h042d191d5a7e1475fc00000000,
104'hb8724c13e4753a8dea00000000,
104'h2c64088fc81665f12c00000000,
104'hbc0b3955163939df7200000000,
104'hb8a16d5a422b0cd95600000000,
104'h30f6c69eed5091f5a100000000,
104'h94e07c0ec01c39493800000000,
104'h28c8e65e91efdf46df00000000,
104'h90b0cff46118231d30a8ece951,
104'hb8367fbf6cdd7c12ba00000000,
104'h9cb9b718731ae5ef3518a50831,
104'h34249aab49d3bc54a700000000,
104'h34703e49e0521d1fa400000000,
104'h60584bd1b05ce9c7b900000000,
104'h940bfd0f17803fc40000000000,
104'h66b3609a6624ffe94900000000,
104'h9486a1b80dbbbcc07700000000,
104'h08a9cb34537d27f3fa00000001,
104'h66323d4f64a5d6aa4b00000000,
104'h2c5bce8db78cf4e41900000000,
104'h90324fa364f53fe0eac770438e,
104'h3480ea4c016d5f77daffffffff,
104'h66e3933ac7f0767ee000000000,
104'h9c0f86e31f2982275309822313,
104'h30fe8966fd33e05f6700000000,
104'h084d61799a611531c200000001,
104'h6600c63301dfa720bf00000000,
104'h28b4b7fa6908aa911100000000,
104'h2c28fc695109541f1200000000,
104'h54da3516b483aa020700000000,
104'h9011c995230d2c731a1ce5e639,
104'h003f9c377f140d012853a938a7,
104'h30b742026e1b4cfb3600000000,
104'h00bf35887e5bdacbb71b105435,
104'h90733cc1e61c8655396fba94df,
104'hb8fbf9f4f76c6459d800000000,
104'h943c5f9978caf8d89500000000,
104'h54027f2d049f406a3e00000000,
104'hbc33eb19679a70a43400000000,
104'h9c06a3970d3507796a04031108,
104'h2c4e468b9ccc81929900000000,
104'h90e9fa62d375cfc1eb9c35a338,
104'h2ca24bfa44cc63429800000000,
104'h00f6f77cedcf693e9ec660bb8b,
104'h60ab543656ae8d0e5d00000000,
104'h34fcdb8cf92d59ad5affffffff,
104'h2c8a02c814701211e000000000,
104'hbcb860027086988a0d00000000,
104'h040fd1ff1f51bd27a300000000,
104'hbc35230b6a5d0b11ba00000000,
104'h30215ee3426aecefd500000000,
104'h3093d38e27aac03e5500000000,
104'h66bb754076502fc1a000000000,
104'h60611d3bc278eccdf100000000,
104'h34a6dba64d699fbbd3ffffffff,
104'hbc69547bd21ca7393900000000,
104'h9ca6df5e4d54feb7a904de1609,
104'h66b4e27c69d563beaa00000000,
104'hb8aea0745d6f9255df00000000,
104'h3419712d3249305b9200000000,
104'h60691db7d263bfefc700000000,
104'h908bd732171ab0c9359167fb22,
104'h902000af4056689fac766830ec,
104'h001ec4013d94da8229b39e8366,
104'h9ccd29aa9a1005432000010200,
104'h545a2bbdb42870c95000000000,
104'h00e2fbb2c53d82777b207e2a40,
104'h04577357ae3740936e00000000,
104'h301768992ea4dc984900000000,
104'h28ce5c789c691c9fd200000000,
104'h043dbce37be97bbed200000000,
104'h54feb190fd86996a0d00000000,
104'h28fb2be0f63c4fcb7800000000,
104'h2c22b1c94595892e2b00000000,
104'h9ce21b9ec413ac572702081604,
104'h54d63d0cacb337e66600000000,
104'h084030e780c6e4be8d00000000,
104'h049ec00a3de86752d000000000,
104'h90ab1b4456a9a81c5302b35805,
104'h047fe02dfff30aece600000000,
104'h9418210530031d4f0600000000,
104'h5448e79f91c1c3ee8300000000,
104'h340a6b3514fcbef0f900000000,
104'h0806f14f0d1d1d593a00000001,
104'h2c24119f4864f75fc900000000,
104'h28c7d4e68fba87e27500000000,
104'h2c25e6d14be17cb4c200000000,
104'h9099d2d433b5160a6a2cc4de59,
104'h042a041554ed6cceda00000000,
104'h30740043e827f80d4f00000000,
104'hb8a515764abf29487e00000000,
104'h0073731de666b7e5cdda2b03b3,
104'h287a65c5f4f1f37ce300000000,
104'h04992e10320f354f1e00000000,
104'h042eaa895d8f488a1e00000000,
104'h54f4cc88e9f161c4e200000000,
104'h340590110bd3fd4aa700000000,
104'h2ce7eeb0cf88bc861100000000,
104'h289605662ccd1a5a9a00000000,
104'h04ee6576dc838e8c0700000000,
104'h9021485742a878165089304112,
104'hb8171e852e93e6942700000000,
104'h04b8b16e71551a9baa00000000,
104'h9c19d0493386551a0c00500800,
104'h2cfe3ff8fccf4dc29e00000000,
104'hb8b565ec6a5a685bb400000000,
104'h940be6011734812b6900000000,
104'h54c32b5c86d8e850b100000000,
104'h34cd94549b7ae42df5ffffffff,
104'h9c2ab94755e3d2b8c722900045,
104'h08da067eb468c1e9d100000001,
104'h94a2a114457c170ff800000000,
104'h54964ecc2c279d374f00000000,
104'h08e9d8f4d339128d7200000001,
104'h2c302249608f0cb41e00000000,
104'h90e5e7cecbadcc305b482bfe90,
104'h54bae4be750356bf0600000000,
104'h34d1d154a3f7f0b8efffffffff,
104'h547b74bbf683cd700700000000,
104'h9469c1edd3748e9de900000000,
104'h342eb78b5d44eaa78900000000,
104'h30bf7ac67e56921bad00000000,
104'h9cd6e53aadf22bfce4d22138a4,
104'h28237dcd469b012e3600000000,
104'h605b9495b773aecde700000000,
104'h544ef9ad9d96f7922d00000000,
104'h0408872511d38c36a700000000,
104'h30ba75d0741b62c73600000000,
104'h90b735366e9ef5123d29c02453,
104'hbccd3e669aea7e04d400000000,
104'h9c2f19d95edf0dfebe0f09d81e,
104'h30519059a3fb0e46f600000000,
104'h9c08bed511858b560b008a5401,
104'h90598553b3c55e4a8a9cdb1939,
104'h2c1f88b93fe90d36d200000000,
104'h6080bfc00195fa8c2b00000000,
104'h545e42cfbcad3b7a5a00000000,
104'h2836d6d16da22d484400000000,
104'h90726b25e432a1bf6540ca9a81,
104'h2c7e826ffd5a3a7bb400000000,
104'hbcb23e82646a4b5dd400000000,
104'h664d87439b355bdf6a00000000,
104'h9441847983a91f745200000000,
104'h287962bdf2f37ceee600000000,
104'h90411b5382d6fcdead97e78d2f,
104'h2cdcb708b910b6eb2100000000,
104'h6695441a2a1596392b00000000,
104'h3421771142e68ccacd00000000,
104'h948eae9c1dbb0dde7600000000,
104'h285bd281b7b6e74e6d00000000,
104'h34824566043c51ed78ffffffff,
104'h5461e1c7c39cd0ee3900000000,
104'hb81bb9c33763383fc600000000,
104'h2c8c120a181ef1e93d00000000,
104'h9cf6cfbcedec5a70d8e44a30c8,
104'h944a513f94dfcc38bf00000000,
104'h60cb6a229668b1ddd100000000,
104'hb8b9fa0a73a7b7984f00000000,
104'h3038567f70fef3a2fd00000000,
104'hb8287fdb50c49d888900000000,
104'h66f8d91ef168ac9bd100000000,
104'h662edadb5d7b7541f600000000,
104'h9c10f90d21471d638e00190100,
104'h94d1b3f8a3077fc10e00000000,
104'h9c3c8c1579abd6565728841451,
104'h00d250dea46343c1c63594a06a,
104'h30ad02c45a711393e200000000,
104'h341c3ffb38d749beae00000000,
104'h66e1f466c3bdd8f27b00000000,
104'h30fbc476f70a97f71500000000,
104'h90286b0750d1ce12a3f9a515f3,
104'h0889023e1210ee652100000001,
104'h080cef7319f4da4ce900000000,
104'h2873ea01e7b2c2c46500000000,
104'h9ccc5534982680c14d04000008,
104'h2c1ce52739eafc90d500000000,
104'h348f46981ee8fc46d1ffffffff,
104'h60a641dc4c567109ac00000000,
104'h9cfc90acf9441b7d8844102c88,
104'hbc6a5f11d4111f252200000000,
104'h9c6e2f3ddcdbdcbeb74a0c3c94,
104'h9002986d053d2ba37a3fb3ce7f,
104'h60d518d0aab6ca286d00000000,
104'h54caf25e952f9d015f00000000,
104'hbc17cab92f1015972000000000,
104'h908e86101dfed776fd705166e0,
104'hbc779501ef5174a5a200000000,
104'h30c8ad6e91eed900dd00000000,
104'hb848a6719110bcad2100000000,
104'h04a6ef264df7355eee00000000,
104'h3408d89b11ad3ece5a00000000,
104'h94b7aaa26f5ed20bbd00000000,
104'h94a13bc442e8e3e2d100000000,
104'h54f1840ee329623f5200000000,
104'h045e62ffbc9908863200000000,
104'h2c7f9059ffd2a2faa500000000,
104'h94eb7012d64b19179600000000,
104'h9c7e412dfc9356f62612402424,
104'hb85bdf8fb778edaff100000000,
104'hbc9510f22a2c02b15800000000,
104'h661014bd20a8e62a5100000000,
104'h9418eedb31f16864e200000000,
104'h6600a5a90195c6242b00000000,
104'h9c236acf4696c40e2d02400e04,
104'h94bc6720783a50fd7400000000,
104'hbccaa17c95f1c76ae300000000,
104'hbc2538af4a5ca5cbb900000000,
104'h0065e84fcbb455f2681a3e4233,
104'h34b790a06ff55b6eeaffffffff,
104'h668b397216d800e6b000000000,
104'h54e8c800d18e5c801c00000000,
104'h94315fd16237433f6e00000000,
104'h9ce8269ad075835feb60021ac0,
104'h9422e31b45907db82000000000,
104'h90ceaefc9d5ef625bd9058d920,
104'h28adb3b65beeb2d0dd00000000,
104'h6009aa7113d342aea600000000,
104'h943b96d5773402c36800000000,
104'h608bf50217853a960a00000000,
104'h663f52617e41e78b8300000000,
104'h30120981246b8f3dd700000000,
104'h28a2990245fb30e4f600000000,
104'h3484cd74093a2db974ffffffff,
104'h54a0b62a411bc04d3700000000,
104'h54471d2b8e975aea2e00000000,
104'h66b9fa0473a204fc4400000000,
104'h04fa17b0f4288f6b5100000000,
104'h542be57b574637f58c00000000,
104'h34042ad308531397a600000000,
104'h041a1639343b57ed7600000000,
104'h66e6df18cd4c5b8b9800000000,
104'hbc53f2aba735e5636b00000000,
104'h602f63d35ed62322ac00000000,
104'h046315ffc6745e93e800000000,
104'h2c8ddb0c1bc249f88400000000,
104'h044e7c219c457b798a00000000,
104'hbc5f658fbe1a6f6d3400000000,
104'hbc3e6db97c4829cf9000000000,
104'h34b6eeea6d874e960effffffff,
104'h94ed2c38da614915c200000000,
104'h08b0b9666153da57a700000001,
104'h90905dc62023268546b37b4366,
104'h949caa12392819455000000000,
104'h9ca739524e22b9194522391044,
104'hb84b54b99657c1bfaf00000000,
104'h54d97286b2769d8fed00000000,
104'h6689c7e6136095e1c100000000,
104'h60d2e5d0a55bd263b700000000,
104'h349818e630f47f86e8ffffffff,
104'h60c8045a90bc33d07800000000,
104'h0826afc54dab6c4a5600000000,
104'h600f00111e12b7d52500000000,
104'h0826534f4c38e98d7100000001,
104'h30f9b7a0f3e96a2ad200000000,
104'hbc76f50fedc180648300000000,
104'h04dc6274b8ed284eda00000000,
104'h60413d5382abd1b25700000000,
104'h60ecfcb8d9531d7ba600000000,
104'hb886d7240d09720f1200000000,
104'h2c67735bce0bfead1700000000,
104'h66357c516a7385d7e700000000,
104'h08229005450106a30200000000,
104'h9cc8c16491f71d26eec0012480,
104'h3481a5240356b1d5adffffffff,
104'h0446a1ab8d6d4fdbda00000000,
104'h906ef9e5dd713a81e21fc3643f,
104'h9c22cb2f455b198db602090d04,
104'h00caf6309536d4a36d01cad402,
104'h5454aabfa934f59d6900000000,
104'h087c0eb7f8cba9f49700000000,
104'h60ac37e458a23b224400000000,
104'h600b70e116c395f68700000000,
104'h2c3180ef631c38ff3800000000,
104'h9c7a6edbf485a1e00b0020c000,
104'h301af6e5350511c90a00000000,
104'hbcbcab92795d40b3ba00000000,
104'h54a679984c1257df2400000000,
104'h300306b306754b25ea00000000,
104'h04e12390c2a7695c4e00000000,
104'h08c348a886b8bbb47100000000,
104'h0829d61d537b8c1df700000001,
104'hbc288e9f51552a9faa00000000,
104'h30fa8548f5a7c9be4f00000000,
104'hbc587681b05b09dfb600000000,
104'h544443df88f88b9cf100000000,
104'h94b90afc72b7a1306f00000000,
104'h006a0f6bd41ef6d13d89063d11,
104'h54236f7d4684ca0e0900000000,
104'h9ca65c384c1e08393c0608380c,
104'hb8af4c2e5e6a6bb9d400000000,
104'h00676157ce0f70731e76d1caec,
104'h6082f9fa058db7261b00000000,
104'h94ee248edc1c2fd73800000000,
104'h00d46e92a84a2319941e91ac3c,
104'h543c466f7844f2838900000000,
104'h3006e85d0db028066000000000,
104'h2c1c8e4139562c51ac00000000,
104'h04915a882285bc2e0b00000000,
104'h94d23610a423f4e14700000000,
104'h6019990333448f8d8900000000,
104'hb8baf6ac75e9a38cd300000000,
104'h9cf04472e05207dba4500452a0,
104'h60efd39edf692b6fd200000000,
104'h34d97648b26cfc99d9ffffffff,
104'h9cb0a734612637654c20272440,
104'h28ce2cb09c0d32ff1a00000000,
104'h2c266e794cd9060cb200000000,
104'h0022769544309a0d615310a2a5,
104'h00c8553690f505beeabd5af57a,
104'h343c5fa178d2467aa400000000,
104'h666f81fddfdf3098be00000000,
104'hb8c79c408f072ec70e00000000,
104'h28e5a214cb3028756000000000,
104'h9011f5a3237ca72df96d528eda,
104'h2c7a358bf41e12f33c00000000,
104'h94fc75b2f8d49da8a900000000,
104'h54ea9b2cd5ea356cd400000000,
104'h00ad53185a1b95f737c8e90f91,
104'h60a8dc8451ee50fcdc00000000,
104'h04ee9d46dd546591a800000000,
104'h344d39e19aa5be804b00000000,
104'h30e5a862cbd5afb6ab00000000,
104'h04be76487cce4a949c00000000,
104'hb88f395c1ef52160ea00000000,
104'h905ce38fb97cd197f920321840,
104'h002c71df583c6d4d7868df2cd0,
104'h903c2e3978c19b9c83fdb5a5fb,
104'h008c7c56182407f948b0844f60,
104'h6637e9976f3878897000000000,
104'h28def7eebd0fa39d1f00000000,
104'h086edbb5dda09bf44100000000,
104'hbc7b2493f6086c351000000000,
104'h9071095de258393db029306052,
104'h66c7cef08f710381e200000000,
104'h662c821b5957df7baf00000000,
104'h902ffc735faf3cfa5e80c08901,
104'hbc64ec3bc909958d1300000000,
104'h04d05744a08799dc0f00000000,
104'h3041d0cb8317b60f2f00000000,
104'h30495a5592a685264d00000000,
104'hb83fa7957f0f8b5d1f00000000,
104'hb8e23d4cc4934f902600000000,
104'h608fa3261f73ab93e700000000,
104'hb8e8a09ad108eb991100000000,
104'h28b23cca649a148c3400000000,
104'hb8f8f968f170697be000000000,
104'h04d8808cb17207e7e400000000,
104'h669bbda237f93332f200000000,
104'h0858193bb00da6fb1b00000000,
104'h00634ff7c68b087c16ee5873dc,
104'hbc3e1c5f7c8b4ee81600000000,
104'h9c76abcfed8dbad21b04aac209,
104'h66cc964699bab4887500000000,
104'h3434d1576942a9758500000000,
104'h086ed5fddd99c0783300000000,
104'h545cf17db92bfd5b5700000000,
104'h2c70794de0852b140a00000000,
104'h54e759eacebda5427b00000000,
104'h348338c406b8d87871ffffffff,
104'h047b210ff65411a9a800000000,
104'h90df73aebe7bf481f7a4872f49,
104'h942c9213592cb0c95900000000,
104'hbc8b7c161614cec92900000000,
104'h94f058e2e0dc2a9eb800000000,
104'h9c15a2cb2b6076abc000228b00,
104'h08ef6e2cde7e5ce7fc00000001,
104'h54cd03549aaa17465400000000,
104'h9ca7c35a4f9c171c3884031808,
104'h2c4510038a1e13753c00000000,
104'h5485ae9a0b82967a0500000000,
104'h2cafddde5ff4e1d2e900000000,
104'h9c6216d5c488c1fe110000d400,
104'h2c5b30b5b631a8bd6300000000,
104'hb8115fbb227e2667fc00000000,
104'h005c4711b8909a4e21ece15fd9,
104'hb8ef15b2de3fb22b7f00000000,
104'h663666416c0110650200000000,
104'h9c1259ed242e31895c02118904,
104'h2808265110c7689a8e00000000,
104'hb8970e522e028a7d0500000000,
104'hbc8b7e0a1622a04b4500000000,
104'h6627c1934f3bb8c17700000000,
104'h00f48efae911b09523063f900c,
104'h9cb45b16682289d54520091440,
104'h607b316df694aa502900000000,
104'h9401870d031f18f33e00000000,
104'hbc1b406f3685921c0b00000000,
104'h607ce25ff9dc0b14b800000000,
104'h54d7a5caafe4fc54c900000000,
104'h9081e6b803738af9e7f26c41e4,
104'h2c8c260e183669156c00000000,
104'h94fb9686f7a2051a4400000000,
104'h6019ec85334860399000000000,
104'hb80ee8f71dbaa3b67500000000,
104'h287ad73bf5844d5c0800000000,
104'h9439f5f573d98ac8b300000000,
104'h000782f90fa21bda44a99ed353,
104'h0813e229278fd40c1f00000000,
104'h9cfc174ef85b92d3b7581242b0,
104'h60998b0233054afd0a00000000,
104'h3407d2890f7b711df600000000,
104'h90b2f2ae654be8d997f91a77f2,
104'h547355b1e6644957c800000000,
104'h345d6c17ba611099c200000000,
104'hb829b09353eb1ddcd600000000,
104'h08a686e64d188afd3100000001,
104'h34b02dbc6021bccb43ffffffff,
104'h0863bb8dc7ed427cda00000000,
104'h54d8de78b16cdbfdd900000000,
104'h9052d731a573bf57e721686642,
104'hb8bbe6d27701f50f0300000000,
104'h600f27c51eea6386d400000000,
104'h9443899987a8e15a5100000000,
104'h940767f10e2366c74600000000,
104'hbc56f455ad5d3601ba00000000,
104'h2c606b21c0c492968900000000,
104'h006fcb55df2b5fd9569b2b2f35,
104'h9c708981e198be2e3110880021,
104'h662675a34c657f81ca00000000,
104'h343fcbff7f6f0a8fde00000000,
104'hb801290b020c05551800000000,
104'h3438d84571c3de6e8700000000,
104'h2891b61a23060d710c00000000,
104'h60f69cc0ed2fa24d5f00000000,
104'h00ae141c5c857bb00a338fcc66,
104'h04dabc9cb5573c65ae00000000,
104'h604fad1d9fb2d7b06500000000,
104'h9cd8bbc4b1da4cb2b4d80880b0,
104'h2c6569e9ca7ce8cbf900000000,
104'h90a1eae6437b28f3f6dac215b5,
104'h90a47e0a4828121f508c6c1518,
104'h2c1e136d3c7c989ff900000000,
104'h2c23f3cf47f96e84f200000000,
104'h08dce382b9f150f6e200000001,
104'h544ef8439d19ac9b3300000000,
104'h08ec1a16d87930f3f200000001,
104'h6079e733f38baabc1700000000,
104'h2c3e72d37ca83d505000000000,
104'h042617274cd2d306a500000000,
104'h008f52241e135c8f26a2aeb344,
104'h2cc0656e80a537544a00000000,
104'h006f3137debed2e47d2e041c5b,
104'hb8668217cdc56d428a00000000,
104'h60e4c9f4c96a7e4fd400000000,
104'hbcfefbe6fde02a2ac000000000,
104'h9ccf030c9ef7d28cefc7020c8e,
104'h28b00c7060099f2d1300000000,
104'hbcf39be8e7e59518cb00000000,
104'h008123fa023695216db7b91b6f,
104'h546698b5cd9d592c3a00000000,
104'h00b3359466cd48a49a807e3900,
104'h94b66e5e6c0ebbc91d00000000,
104'h601bc309372a06155400000000,
104'h0808ee9311d45fa4a800000000,
104'h348ea8e41db3858c67ffffffff,
104'hbc14f3b929dea93ebd00000000,
104'h0022aa7345db06e8b6fdb15bfb,
104'h2ca4cd0049603ad3c000000000,
104'h28dcbdbeb9242dc34800000000,
104'h660d6a551a78305df000000000,
104'h540e17971c109d7b2100000000,
104'h00c648628cd61b98ac9c63fb38,
104'h0470f785e18b55281600000000,
104'h300e1c951c53c001a700000000,
104'h34d033d6a02fcbad5fffffffff,
104'h3448411990408ed58100000000,
104'h00c585968b88cb9e114e51349c,
104'h087ee0d7fddae30cb500000000,
104'h00da9490b5230f5d46fda3edfb,
104'h0035e3816b32fd676568e0e8d0,
104'h2c18c353310f9d031f00000000,
104'h667a997df573c05fe700000000,
104'h94d3bb26a731e26d6300000000,
104'h28dc27fab84d2c319a00000000,
104'h943ab81975759135eb00000000,
104'h34b8b4e671fc9ad8f9ffffffff,
104'h08fc94f6f9c83aba9000000000,
104'hbc0b52e9162ebc135d00000000,
104'h9c0a974b1572ac17e502840305,
104'h04a6ad704db7515a6e00000000,
104'h2845fb618b2e0a295c00000000,
104'h2c8874aa10daa9eab500000000,
104'h04a440464810ad892100000000,
104'h08b1898063a4dec24900000000,
104'h301633c92c2ebe955d00000000,
104'h90aee99e5d8ace9a1524270448,
104'h903dbe6f7b8a916815b72f076e,
104'h28bf5b707e50d9f1a100000000,
104'h04be6f887cb0c1e06100000000,
104'h0041da2583f35f00e635392669,
104'h54b4c922691c0f973800000000,
104'h2cd8c1a6b10cf5c71900000000,
104'h28a04c04403cf9eb7900000000,
104'h346dba9fdbf66bfcec00000000,
104'h9ccc43c098c11bf482c003c080,
104'h9402667f049c81223900000000,
104'h9c03529d06764895ec02409504,
104'h54f9cb6cf3c762728e00000000,
104'h9419bda933e56662ca00000000,
104'h544680598d4fe6e79f00000000,
104'h669a78ae34810bbc0200000000,
104'h04a998ec537e8b3dfd00000000,
104'h94a2f23c4503dabf0700000000,
104'h60ee5196dc902df02000000000,
104'h2cb99f9c735a9d45b500000000,
104'h54ce7b809c1c8b3f3900000000,
104'h602b48db563620e96c00000000,
104'h54eba896d7da7922b400000000,
104'h2c3b14c57620d30b4100000000,
104'h9409178712fde358fb00000000,
104'h083154e562b41cc26800000000,
104'h04725fbbe42b875d5700000000,
104'h301511892a497ef19200000000,
104'hb83add5f75be70687c00000000,
104'h669c55ba38436e2d8600000000,
104'h9cc1dd6083db337ab6c1116082,
104'h089f3b463ec9eed49300000001,
104'h66a7896a4f8ceb501900000000,
104'h9c19b6bb3396f1042d10b00021,
104'h081e93eb3de7f462cf00000000,
104'h34882360102e6c995cffffffff,
104'hb846a40b8dee68eedc00000000,
104'h042a8f45559e3d2a3c00000000,
104'h08fb81b6f7b25cf06400000000,
104'h287ac735f5a1be1a4300000000,
104'h3445019d8af1da22e300000000,
104'h60e122bac2c526808a00000000,
104'h0453b127a7289c055100000000,
104'h04741025e8e4a53cc900000000,
104'h94b642806cd38bcea700000000,
104'h904e607b9c233ce7466d5c9cda,
104'h3433b8996761fc81c300000000,
104'h66c8538e90355fdd6a00000000,
104'h60765319ec10a6d32100000000,
104'h949f63e63e9b4c3a3600000000,
104'h9c733a6fe6aa65425422204244,
104'h28d8d2d2b12727db4e00000000,
104'hbc3aebc575eab00cd500000000,
104'h30eaf45ed5eadc5cd500000000,
104'h9c9e65063cfdd92cfb9c410438,
104'h00793b55f269b31bd3e2ee71c5,
104'h2cd510e2aa5b085fb600000000,
104'h60af05405ea9b12e5300000000,
104'h900f72c31ef3f71ce7fc85dff9,
104'h0005266f0a80b3760185d9e50b,
104'h94a292d445766ca7ec00000000,
104'h54fe35ecfc394a917200000000,
104'h54382a01701b79f53600000000,
104'h082599854b6b56d5d600000001,
104'h942f8df95f4075c78000000000,
104'h665d51c5baa464604800000000,
104'h301b5d2336c5b8948b00000000,
104'h604685f78d3bc70f7700000000,
104'h0807eaaf0fef189cde00000000,
104'h0450d027a16e767fdc00000000,
104'h54f66a88ec4225db8400000000,
104'h54bc4922789eaa0a3d00000000,
104'h00b8dd58719e26083c570360ad,
104'h2c9a5474345334cda600000000,
104'h601abc8f3589d0a61300000000,
104'h9c992c6a3252a1a3a510202220,
104'h540266570472caede500000000,
104'hb8262e0f4cf60f2aec00000000,
104'hbcf7499aee5ae3dbb500000000,
104'hb832e52d658fcbbc1f00000000,
104'h0438d207712f10295e00000000,
104'h90a8d8525181b1760329692452,
104'h66521407a4c426548800000000,
104'h905814cbb05f4233be0756f80e,
104'hb8d638c8ac355a9b6a00000000,
104'h66ec7aa0d83783916f00000000,
104'h94b1aa3863207af74000000000,
104'h2c35c8a36be29aeac500000000,
104'h603bfeff77fbeb24f700000000,
104'h28ce685a9cef295ade00000000,
104'h2cf6a68ced82609e0400000000,
104'h2cecfa16d98b67be1600000000,
104'h94a4550848f05ea4e000000000,
104'h00eca0ded98602b20c72a390e5,
104'h34252f634a8f722e1e00000000,
104'h66d80e84b042b6958500000000,
104'h9443b74587cb2dfa9600000000,
104'h54034f8f063eab7b7d00000000,
104'h285e771dbccbe6869700000000,
104'hbc80574c008091460100000000,
104'h669a6e1434532e0ba600000000,
104'h60fa4bcaf4107b932000000000,
104'hbc0a3c1914561083ac00000000,
104'h044391d387537dbba600000000,
104'h94f60dd6ec910fae2200000000,
104'h08a298f045e706d8ce00000001,
104'h343048b96011df092300000000,
104'h90a967705257fdcbaffe9abbfd,
104'h6622f6eb4572dfcbe500000000,
104'h2c23e66147d19d2ca300000000,
104'h2801f35b03445cf58800000000,
104'h0868ed8bd1a00f5a4000000000,
104'h9c4dd5b39bdf873ebf4d85329b,
104'h341a0f7d3422ca714500000000,
104'h90939e60279f31263e0caf4619,
104'h301e25813c8aac4a1500000000,
104'hbc15228f2a3a4ae97400000000,
104'h28629ba3c57fd685ff00000000,
104'h30c638288cbc1e807800000000,
104'h2caf7cb05e8b4a781600000000,
104'h08caa1dc95564babac00000001,
104'h349a3e3434e04546c0ffffffff,
104'h6060bb15c10883e11100000000,
104'h04634c7dc6e15bc6c200000000,
104'h54e4e3fcc9da0662b400000000,
104'h2c4a5693947d5697fa00000000,
104'hbc59ad83b320dc294100000000,
104'h28a55a424a3fce137f00000000,
104'h00a0c5504112d3f125b3994166,
104'h94c6701a8cb186566300000000,
104'h0850a1d5a19c3e363800000000,
104'h007c5765f8648b3fc9e0e2a5c1,
104'h08d2ee38a53869377000000001,
104'h60b9c22c73c80c669000000000,
104'hb837b6696f47dced8f00000000,
104'h34af61405e9ff9283fffffffff,
104'h30e95312d22057154000000000,
104'h3064b02bc9bc5ca47800000000,
104'h902d15a15ad2872aa5ff928bff,
104'h669b8138374c79b39800000000,
104'h901cb44139618a69c37d3e28fa,
104'h9c8a497414e9a6f0d388007010,
104'hb88475da08e827ccd000000000,
104'h94b92caa7235eabb6b00000000,
104'hbcd21e20a4e7cc14cf00000000,
104'h540dc9671baa572c5400000000,
104'h3400997901bd45b87a00000000,
104'h66d1c4f6a3f12622e200000000,
104'h602c691358f740f6ee00000000,
104'h9440176780e79538cf00000000,
104'h283cced9790a83cb1500000000,
104'h90e51780ca2381c947c696498d,
104'h30cdb9789b9fe9ee3f00000000,
104'h34dd46d0ba98c4f231ffffffff,
104'h9046705d8c7820e3f03e50be7c,
104'h66bedda27dba4f8e7400000000,
104'hb8c8ffb291a123e04200000000,
104'h04ba17047433063b6600000000,
104'h00666465cc7977e3f2dfdc49be,
104'h903c3cc178125d53242e61925c,
104'h90c3781e86bd27a67a7e5fb8fc,
104'hbc2173654208b4f31100000000,
104'hbc1a9d4d35987fa83000000000,
104'h9c41463b820f74f71e01443302,
104'h94462b1d8c7c8a25f900000000,
104'hb8e1f350c398e8fa3100000000,
104'h603f997b7f314b176200000000,
104'h2c5e776fbc23dc594700000000,
104'h343f6d0f7e61bc3bc300000000,
104'h9c0b5a2516cef6309d0a522014,
104'h2c69e349d39d890a3b00000000,
104'h082639bf4c47d55b8f00000001,
104'h60b45e54688c8ac61900000000,
104'h9c5c1747b831ec756310044520,
104'hbc6f911ddfd00466a000000000,
104'h0432628964e11ddac200000000,
104'h00a26b4c44cd9eaa9b7009f6df,
104'h2c5ec613bd0417a90800000000,
104'h9421c5534360240bc000000000,
104'h66d9b32eb39a6fba3400000000,
104'h2c10cc572129fcc55300000000,
104'h0837ade96f527fada400000001,
104'h94362e4b6c056ad50a00000000,
104'h9095590e2a2b00d956be59d77c,
104'h345205d7a4ce85f49d00000000,
104'h0022422b44f4685ee816aa8a2c,
104'hb8608667c182f7a40500000000,
104'h90166d8b2c0e03171c186e9c30,
104'hbc756827ea73771de600000000,
104'hbc9ea2383d7ad19ff500000000,
104'h2c9c14043803055d0600000000,
104'h2c0b7601162a24535400000000,
104'h30e88faad12fe91d5f00000000,
104'h284f19719e0ff74f1f00000000,
104'h54a529864ae26adac400000000,
104'hbc95e3d22b690e6fd200000000,
104'h0048e4c391bd50d27a0635960b,
104'h90859f320b46d14f8dc34e7d86,
104'h08a2a54a45ec1b00d800000001,
104'h606f945fdf3ee7497d00000000,
104'h30651bcdca2aff215500000000,
104'h9c8156e002da937cb580126000,
104'h00ff71b2fe04a4ad0904166007,
104'h04c051048021d0c34300000000,
104'h346eb529dd01a0e50300000000,
104'h005c0fd9b85e2db9bcba3d9374,
104'h5474051de845b2c18b00000000,
104'h66a34f2846f168bae200000000,
104'h005b7d39b6d6befead323c3863,
104'hbca7c57c4fdbcbe4b700000000,
104'hbc3fe1eb7f898c1c1300000000,
104'h2c5cb025b94e49139c00000000,
104'hbc770c5dee503e53a000000000,
104'h00bc1f2c786455e1c820750e40,
104'h9493167a2666939dcd00000000,
104'h083f015d7ee187a8c300000000,
104'h9c2446f34897dfba2f0446b208,
104'h28b3f046678eef8a1d00000000,
104'h2827bd2f4f9ac8263500000000,
104'h6640bc318194365e2800000000,
104'h34cedd5a9d3ec01b7dffffffff,
104'h901ab82b35e878c2d0f2c0e9e5,
104'h900b7c6516e74496ceec38f3d8,
104'h0841c5ff83b6e3126d00000000,
104'h280ccbf91990d8522100000000,
104'h044a223b94530d6ba600000000,
104'h2899067e325bbfcdb700000000,
104'h0000f029011917a7321a07d033,
104'h90efdb26df587d41b0b7a6676f,
104'h607785d5ef558561ab00000000,
104'h60a199da43120cab2400000000,
104'h00c1780c8210d9f921d25205a3,
104'h66871f480e11dfc72300000000,
104'h3071665be25af487b500000000,
104'hbcc680da8d599a0fb300000000,
104'hbca0870c41722bebe400000000,
104'hb89078be208e8cc21d00000000,
104'hbc0cf32d19e22abcc400000000,
104'h540291dd0552f2dba500000000,
104'hbc9ab28635768b5bed00000000,
104'h285a13e7b408ed151100000000,
104'h944387a9879d33e03a00000000,
104'h5463af43c7fb3decf600000000,
104'h28417bdd8294722a2800000000,
104'h94d3e920a7a7c59e4f00000000,
104'h28002b2f0080d7d20100000000,
104'h60f4476ce8a7be264f00000000,
104'h5420d06d4146d6398d00000000,
104'hb8d13ccea271b741e300000000,
104'h609d11203ac41a748800000000,
104'h08d4d4b6a9f15268e200000001,
104'h00d48996a9c4a966899932fd32,
104'hb87a1f51f4b0bed86100000000,
104'h901118dd22cfbba69fdea37bbd,
104'h66855d860a0ff5911f00000000,
104'h66cdecbe9ba859925000000000,
104'h04eced04d9c5b5488b00000000,
104'hbccd4dc49a1db7473b00000000,
104'h085ef437bda63e7e4c00000000,
104'h60c92b3e9287509e0e00000000,
104'h900fce4b1f6bcf6fd7640124c8,
104'h304a67399408c5351100000000,
104'h043d372d7afce014f900000000,
104'h94f2e27ae5797469f200000000,
104'h54923784246c1e2bd800000000,
104'h2c4648978c8bd9521700000000,
104'hbc57d0c5afae29305c00000000,
104'h00bd9bd27b90a6d2214e42a49c,
104'h281e69133cc10e608200000000,
104'h08b1813e63f1a380e300000001,
104'h664bf75f97c184b48300000000,
104'h08674ca5ce4045bb8000000000,
104'h2cbaef527529e8eb5300000000,
104'h604ccc9399740f9de800000000,
104'h0455ed5dab36f97f6d00000000,
104'hbc2ed6535db4ab026900000000,
104'h345c22a7b82e52ad5c00000000,
104'h60f691f0edcbc5869700000000,
104'h9cba811c7502aa710502801005,
104'h0839863b731aac893500000000,
104'h28a5a76c4b91cc862300000000,
104'h04a864ba50afa9205f00000000,
104'h08608d01c178566bf000000001,
104'hb82895bf51d71c2eae00000000,
104'h30dbee04b73733576e00000000,
104'hbc24845149445a4b8800000000,
104'h2c9a77663426d8494d00000000,
104'h045eaa3dbdae47d25c00000000,
104'h6005b2d10b743fffe800000000,
104'h34535c11a67bb4e3f700000000,
104'h9c1fb2b13f23a6f14703a2b107,
104'hb8f55516eadb7956b600000000,
104'h9c3d7e317ad5075caa1506102a,
104'hb851035ba26450c9c800000000,
104'hbc363d3d6cc6553e8c00000000,
104'hb86293abc51876993000000000,
104'h60332483664f7a519e00000000,
104'h082abd91556901dfd200000001,
104'hbc0c216d18d41212a800000000,
104'h28ce4f5a9c95017a2a00000000,
104'h9cdd4626bae6e5bccdc4442488,
104'h944c7a11988058040000000000,
104'h0440f59f811b284f3600000000,
104'hbc17dd852fde57dabc00000000,
104'h305acf7fb5bf72807e00000000,
104'h009e543c3c4c1f1998ea7355d4,
104'hbc9f5c343e7e7ed1fc00000000,
104'h2c8b7f8816b6b3986d00000000,
104'h280478eb08a1a57a4300000000,
104'h54521375a428defb5100000000,
104'h9006838d0d71187be2779bf6ef,
104'h2c47e2cb8fdcca98b900000000,
104'h9cae46c85ceddf8cdbac468858,
104'h6060ab17c12d5b8d5a00000000,
104'h3483a60807e1942ac3ffffffff,
104'hb853a0a5a7c34eb48600000000,
104'h6019097b32ffdd94ff00000000,
104'h66b7ba826f1a14af3400000000,
104'h2c9b8a063795acc22b00000000,
104'h3062be7bc5386dd37000000000,
104'hb893dd5e270238750400000000,
104'h2c170d1b2e38c63f7100000000,
104'h2cc401e888f5b922eb00000000,
104'h9c4c2dad98fd51ccfa4c018c98,
104'hb8cdaad49b31e50b6300000000,
104'h9c9e1a3c3c2be81d570a081c14,
104'h000d6c0f1a482c2990559838aa,
104'h542f4b995e4da0899b00000000,
104'h00d6a63ead91b43623685a74d0,
104'h0809854b13ae2e2a5c00000000,
104'h54fc32d4f85d14b5ba00000000,
104'h604961a19256fbe1ad00000000,
104'h3451cffda30dd2db1b00000000,
104'h9ca09da4414208498400080000,
104'h9c924ca024a99da853800ca000,
104'h607b2523f6a081ba4100000000,
104'h08d6746cac0f49d71e00000001,
104'h94d2dea8a5d12254a200000000,
104'h0488bbcc11d38de2a700000000,
104'h607e3781fc624bf1c400000000,
104'h0081abee037f7e09fe0129f801,
104'h30856fb60a3be42f7700000000,
104'h60b90ebe72acc8445900000000,
104'h94caa61895ccf0689900000000,
104'h08b7dae46f3bb0537700000001,
104'hbc10a43121d8f1b8b100000000,
104'h94b6dfd26d9ecbac3d00000000,
104'h662c6a4d584100fd8200000000,
104'h9c1631af2cf87d92f010318220,
104'h90ed7b74dae4aad0c909d1a413,
104'hbc995568328632fc0c00000000,
104'h3408e97b11768b93ed00000000,
104'h90942caa28955ea82a01720202,
104'h341320e526e0ab58c100000000,
104'h34f4a1e2e9fe3514fcffffffff,
104'h04547503a8949a042900000000,
104'h08d5143aaae02878c000000001,
104'h54046be108e34b30c600000000,
104'h0003839f071c24d1381fa8703f,
104'h9437ca496f38b2397100000000,
104'h90a97cbc52c88bdc9161f760c3,
104'h9c8d5fc61ad71e36ae851e060a,
104'h3000c4ff019af1163500000000,
104'h046592a7cb6e5609dc00000000,
104'h30c0c690810395b90700000000,
104'h6630abf761aa744a5400000000,
104'h30b0bc606176a4c3ed00000000,
104'h341fe3813f9683582d00000000,
104'h548a9e18151f2eed3e00000000,
104'h00452bd38a6ed94fddb4052367,
104'h601acc2735f7e6b4ef00000000,
104'h28edbe36db3f34097e00000000,
104'h04487bb590059c570b00000000,
104'h34c366b886689523d1ffffffff,
104'h3072e2afe52f79cf5e00000000,
104'h5400902701eaddf6d500000000,
104'h284f23c39ef0fed8e100000000,
104'h30c3100a860e2ba51c00000000,
104'h0432fa5b65e1bceec300000000,
104'h0449b2b393c7f3048f00000000,
104'h907826a3f0ced3509db6f5f36d,
104'h2ca8872851f7dcb4ef00000000,
104'h9c649989c9e22af6c4600880c0,
104'h903feb397f586111b0678a28cf,
104'h54c360b68613729f2600000000,
104'h0802577104bf24347e00000000,
104'hb81a529b34dedac4bd00000000,
104'h9c54eb1ba90911fd1200011900,
104'h08287a5f50fd91a4fb00000000,
104'h3416b8432dce3a049c00000000,
104'h941943ef329bff3a3700000000,
104'h041acfb735b96ba67200000000,
104'h609867f83049c1439300000000,
104'h30210d01421f92033f00000000,
104'h9cb297e6659f67383e92072024,
104'h6019a26f3332cff16500000000,
104'h002ee9e75d55ee57ab84d83f08,
104'h083f650b7eed5c0eda00000000,
104'h30cd04e09a4bfd9b9700000000,
104'h9c54d8a1a9901cb8201018a020,
104'hb8940c8628b4e1c26900000000,
104'h660ffbbd1f51040ba200000000,
104'h001e4d3f3c6d4947da8b968716,
104'h9c80d3ac01952be02a8003a000,
104'h288da8381b31c0656300000000,
104'h08feb87cfdd2b1d6a500000000,
104'hb894bf5e2932ed196500000000,
104'hb8e860f6d0f65346ec00000000,
104'h9cc0e15e81438b1d8740811c81,
104'h6042aea785e8c950d100000000,
104'h66f0b5a2e19c27f03800000000,
104'h000239d9048fe4cc1f921ea523,
104'h2ca3a85847f09ecee100000000,
104'h668b9d9a17676a59ce00000000,
104'h9c8e166a1c5354b1a602142004,
104'h30b683b66d8dae501b00000000,
104'h049e39843c2234554400000000,
104'h285f70bbbedff0d0bf00000000,
104'h085dd413bbf96a36f200000000,
104'h08544ff1a88279b40400000000,
104'h045c9d43b967e093cf00000000,
104'h9c27bf674ff07498e020340040,
104'h540f6d011ee17b64c200000000,
104'hb8371be56e6f8cd7df00000000,
104'h9c5027f5a02b14695600046100,
104'h30ef4cfade83498e0600000000,
104'h2c6a6b8fd43c37197800000000,
104'h601c50f538bc29987800000000,
104'h3060f9fbc1529cb5a500000000,
104'h54cf88dc9ffe7f92fc00000000,
104'h04d7e622afb368346600000000,
104'h9428c47f511d0dd93a00000000,
104'hb8cf7fb29e562259ac00000000,
104'h040e0e691c636287c600000000,
104'h9c1bff1937757599ea11751922,
104'h089e37e43c6bf379d700000001,
104'hbc45f17d8bc1aa328300000000,
104'h04ea24fed45dfa4bbb00000000,
104'h043f64d17eb0e2226100000000,
104'h9040d885816f1057de2fc8d25f,
104'hb819d3bd332915235200000000,
104'h661a400134448abd8900000000,
104'h28a8d1ac517fccb3ff00000000,
104'h9c6cbfc1d99096542100964001,
104'h60bd76cc7a8ba00a1700000000,
104'h00f97ecef20713bd0e00928c00,
104'h34668c0bcd43702b8600000000,
104'hb8db72f6b68633500c00000000,
104'h66617711c22763cb4e00000000,
104'h90652cc7ca0ed12d1d6bfdead7,
104'h60a7e64c4f6fa369df00000000,
104'h3019638932e8912cd100000000,
104'h30c63ce88cbcd5407900000000,
104'h944a4149940dbaed1b00000000,
104'h2c66bed1cdc6594e8c00000000,
104'h90ab6ed456bad5c67511bb1223,
104'h003d7cb37a42454f847fc202fe,
104'h30e2dfb6c5be04da7c00000000,
104'h6640fff9810320bb0600000000,
104'h34e45e3ac8e22300c4ffffffff,
104'h90dbb6ceb70760d30edcd61db9,
104'h66a3d76e47919ed62300000000,
104'h0082202204f6a48eed78c4b0f1,
104'h2c6a671fd48d16b81a00000000,
104'h60d9b79eb348b0ad9100000000,
104'h66da23d2b451b4c3a300000000,
104'h085ca1b1b9122bab2400000000,
104'h046caadbd98b4ad01600000000,
104'h602617834c3319c16600000000,
104'h66f86c42f0ae2e7e5c00000000,
104'h04539301a76318ebc600000000,
104'h6088b6d21194d5262900000000,
104'h0426bad94d575ce9ae00000000,
104'h0094841c29bd2fe87a51b404a3,
104'h08d40e74a8fe6b34fc00000001,
104'h34600467c081c79c0300000000,
104'h34aa5200548d97081bffffffff,
104'h5414eac1296a98e1d500000000,
104'h34feba6afddc3d64b8ffffffff,
104'h04dd78f4ba71b011e300000000,
104'h2809d95f1348c1019100000000,
104'h900e4b911cd78548afd9ced9b3,
104'h9ca149444223465b4621404042,
104'h302ae5df55e31864c600000000,
104'h667a194df45a2fafb400000000,
104'h0450fdeba1a9ccfe5300000000,
104'hbc5ff961bfe458f8c800000000,
104'h28568883adbb06767600000000,
104'h9c8d262e1a2513f54a0502240a,
104'h90a685304d4b83e597ed06d5da,
104'h2c0f15211e45e41d8b00000000,
104'h00a88a42513c7c2978e5066bc9,
104'h34e3e064c741fab183ffffffff,
104'h543f10c37e1a79db3400000000,
104'h543c72e3781f72a93e00000000,
104'h04a8807c51eff758df00000000,
104'h000f744d1e924cc224a1c10f42,
104'h94cefbfe9d87babe0f00000000,
104'h00e8f508d1052b7b0aee2083db,
104'h34d2ec92a57af1e9f5ffffffff,
104'h90a2da4645c3cf0c8761154ac2,
104'h945c4e45b8270e714e00000000,
104'h947209f3e4c351748600000000,
104'h94febbe2fd6761b7ce00000000,
104'h667456b5e844226f8800000000,
104'h90bc3af678ae78d25c12422424,
104'h28ab2bfc5649c3779300000000,
104'h0072c7cde5db38a4b64e00729b,
104'hbc0ef9f71da443c64800000000,
104'h94c0a17281e5b9c4cb00000000,
104'h0027618d4e077c5f0e2eddec5c,
104'h90ab55b4563fe4917f94b12529,
104'h0454206ba86c0bf7d800000000,
104'h08158d1b2b85cd240b00000000,
104'h2cb2bcfc65b6130c6c00000000,
104'h2ccf96f49fd9cf5cb300000000,
104'h044cf271995dafddbb00000000,
104'h66ceb54e9d086ad31000000000,
104'h30fbdcb2f7953a622a00000000,
104'h60d728f0ae4fdee79f00000000,
104'h662be46b572940595200000000,
104'hb8a4fd6c496786b1cf00000000,
104'hbc6d6b0bda16413f2c00000000,
104'h905f9509bf22f511457d6018fa,
104'h667e36b9fc902a4e2000000000,
104'h04e3f4d4c7ccd09e9900000000,
104'h90379e656ff79282efc00ce780,
104'h9431d09b63156fb92a00000000,
104'h9c8d75b81af8b698f188349810,
104'h900756e90e31347b623662926c,
104'h2c89b92213d0350ca000000000,
104'hb877bd09ef82a8c00500000000,
104'h04f0f9cce1718a1be300000000,
104'h30088b0711ec5a24d800000000,
104'h34fb89a2f70b4bbf16ffffffff,
104'h90a1a7b043a676064c07d1b60f,
104'h344f67539e2525b54a00000000,
104'h605c2491b834257f6800000000,
104'h6626ea474d539579a700000000,
104'h00fbc9f4f7d4a96ca9d07361a0,
104'h08502eaba03d66457a00000000,
104'h549f62e63e8c36681800000000,
104'h9471416de26eed17dd00000000,
104'h30f3c932e7a090d04100000000,
104'h66bd0c367a3704ad6e00000000,
104'h2cf5b166eb2568c14a00000000,
104'h080501770a89c97e1300000000,
104'hbc0e36cd1cf47614e800000000,
104'h2cd38856a7a515ca4a00000000,
104'h041627712c2d54675a00000000,
104'hb8fb28c2f6f2bd8ce500000000,
104'h908c102018191f1732950f372a,
104'hb8c677688c648a7fc900000000,
104'h04090867120dcd3d1b00000000,
104'h9cb4c1b26945f8218b04c02009,
104'h30c03e9080ad4db85a00000000,
104'h666f79cdde3fafab7f00000000,
104'h609543a62a9c63223800000000,
104'h306462a5c808c41d1100000000,
104'h3015177b2a8d3fd81a00000000,
104'h60307be56001ae2f0300000000,
104'h045df493bb39e1f77300000000,
104'h08c7adfa8fb5085e6a00000000,
104'h60c1dc3e83aa2f565400000000,
104'h080536110afa0ae8f400000000,
104'h94afe28a5fe1d198c300000000,
104'h9010d2132134c7c9692415da48,
104'h94303a4160d1d216a300000000,
104'h9cc4acae89f026bae0c024aa80,
104'h30ff00ecfe29f5eb5300000000,
104'h6000094f00cda1389b00000000,
104'h3411cadb2365d9f3cb00000000,
104'h0092b0202586be820d196ea232,
104'h6613ef192731cecd6300000000,
104'h302d1a0d5a7c4f91f800000000,
104'h342593714b0374d10600000000,
104'h9c815cc4020f6b231e01480002,
104'h2ce97870d282181c0400000000,
104'h9c80d6ae01c029b0808000a000,
104'h30ad85625b1acc8b3500000000,
104'h28629afbc5ce21789c00000000,
104'h003a145374dc49bab8165e0e2c,
104'h08de9d94bdd6a276ad00000000,
104'h2c93fe0e27768707ed00000000,
104'h60c99f2493acb2645900000000,
104'hb8bd66207afa1788f400000000,
104'h08fdd91afb66c8c3cd00000001,
104'hb84146d782b3461e6600000000,
104'h003c69a3785e4ac9bc9ab46d34,
104'h6615bd3b2b3cf1677900000000,
104'h28737fa7e69cc7763900000000,
104'h0021151942a727b84ec83cd190,
104'h549546d22af2f384e500000000,
104'h946d94ffdb4d83339b00000000,
104'hbceb9392d7b565706a00000000,
104'h28d80a36b0b945ae7200000000,
104'h34944f1428db1176b6ffffffff,
104'h08c514cc8aab34cc5600000000,
104'hbc92a34425f98592f300000000,
104'h0829338f522935e75200000001,
104'hbca0e6ca415ae581b500000000,
104'h08ef9006df2baa175700000001,
104'h54af49185e29a6bb5300000000,
104'h548b8a8217468a3b8d00000000,
104'h28bb3e54766e0c81dc00000000,
104'h0441060b826a42efd400000000,
104'h286bab6fd75963cbb200000000,
104'h906f7471de98509030f724e1ee,
104'h549dd2103b1aff573500000000,
104'h90eba23ad7279b374fcc390d98,
104'h34cefca89d3af3a375ffffffff,
104'h663442b968f492c2e900000000,
104'h940eea611d3692e76d00000000,
104'h2c0d3bf71a990ace3200000000,
104'h66e6fb24cddaa91eb500000000,
104'h2ccdb2be9b87d6b60f00000000,
104'h90621ba3c497780a2ef563a9ea,
104'h2c6cd69dd9a825945000000000,
104'h2c21714542ca73249400000000,
104'h66196ddd32cc9e469900000000,
104'h2c29c63753b9bba67300000000,
104'h60e8218cd0223b694400000000,
104'h54d5b566abbd5c907a00000000,
104'h2ce48976c972e757e500000000,
104'h2c18967f31d2469aa400000000,
104'h9490f82821d7d82caf00000000,
104'h60fe29ecfc930c422600000000,
104'h94a106ec4237abc76f00000000,
104'h301304db26525dc5a400000000,
104'h907ae1cff5ac43c058d6a20fad,
104'h5421bd3543d3451ca600000000,
104'h34cb539c96ac617458ffffffff,
104'h0870d5a9e1db2206b600000000,
104'h003891e1719502022acd93e39b,
104'h9c6d69a1da9965fc320961a012,
104'h2cffc8e8ffee7a42dc00000000,
104'h2c6e9949dda1103e4200000000,
104'h080967bf128952d21200000000,
104'h66fdb58efbefe9c4df00000000,
104'h54c02c2e804ee40f9d00000000,
104'h54cf2c1c9e3f814d7f00000000,
104'h54b6eec66d61b213c300000000,
104'h30583361b09be7523700000000,
104'h04e92ed0d2e988bad300000000,
104'h54ad36845afc2a12f800000000,
104'h30225e5944a757a24e00000000,
104'h901501752a589189b14d90fc9b,
104'h34d7ee2caf2cce2559ffffffff,
104'h287cacdff97a9b71f500000000,
104'h008219d60453b761a7d5d137ab,
104'h9cb84a2c7082b7460580020400,
104'h9c3f73a57e51162fa211122522,
104'h9c3c4f8d78dfc244bf1c420438,
104'h344f30a19e80012c0000000000,
104'h60bbc3e6773443696800000000,
104'h9cae34965cc03eb68080349600,
104'h60d72aecae656771ca00000000,
104'hbce2de12c504a0e90900000000,
104'h54c8310490cfbcd49f00000000,
104'h9cc39262876d219fda41000282,
104'hb8b6175e6c5dafd3bb00000000,
104'h28c409928808be751100000000,
104'h081edfe53dfbc666f700000000,
104'h08155a6d2a1b14c53600000001,
104'h9081394402a69c4a4d27a50e4f,
104'hb8a4c67c4981bdae0300000000,
104'hb8332ae9660e9eff1d00000000,
104'h08c5460e8a956a0a2a00000000,
104'h341180ff238d89bc1b00000000,
104'h600fd4311fa2be764500000000,
104'h3473f871e7e9a17ed300000000,
104'h66c67aac8cd6ef4ead00000000,
104'hb8922aea2422b1034500000000,
104'h90c61e108c3c1caf78fa02bff4,
104'h66453ad98a44c4c58900000000,
104'h08d309a6a6216e734200000001,
104'h04d23f68a4fca700f900000000,
104'h00cc3b7c980af03715d72bb3ad,
104'h04297087526a1bb3d400000000,
104'h6011705b22052d550a00000000,
104'h94c612da8c6bdc97d700000000,
104'h3427efd14ff88cecf100000000,
104'h941b23d536615527c200000000,
104'hbc6a182bd4586dd7b000000000,
104'h3438c5a1711e1ea33c00000000,
104'h2c4daa739b4a02b19400000000,
104'h9c166b292c8b3c021602280004,
104'hb88cd674191eedd73d00000000,
104'h9cadc4185b3216076420040040,
104'hbc3e06bf7cbf9d647f00000000,
104'h90d268dea4ad37265a7f5ff8fe,
104'hbca66c9a4c616737c200000000,
104'h9c7246a3e4bac7a0753246a064,
104'h08534c15a6a464e84800000000,
104'h28aacb56556cc971d900000000,
104'h9cc607fa8cf50fd4eac407d088,
104'h2cded1a2bdb314506600000000,
104'h66beedd67dcd9d1a9b00000000,
104'h60b94cf2723b11c17600000000,
104'h28f2c1f6e53319936600000000,
104'h9cc8b572916138f9c240307080,
104'h54b70b646e8a45da1400000000,
104'h2c1f34113eb04af86000000000,
104'hb8f11fece2a0324e4000000000,
104'h66238e77472a4e795400000000,
104'h3453f01da7829b0a0500000000,
104'h607ed313fd574bf7ae00000000,
104'h54b8933e718403ea0800000000,
104'h9cd2c50ea5d5c9aeabd0c10ea1,
104'h2c1d935f3b87948a0f00000000,
104'h90a508564ae9079cd24c0fca98,
104'h3498f94a3170b445e1ffffffff,
104'h60ab0d985640fb7d8100000000,
104'h3449188d92526639a400000000,
104'h0462be3fc5f80cc8f000000000,
104'h2c101b7120ba653e7400000000,
104'h60a3e874478290c00500000000,
104'h04a64f044c33fff56700000000,
104'h04966b282c0c065d1800000000,
104'h004f2f159edeb4b6bd2de3cc5b,
104'h08392205727e125bfc00000001,
104'h9c3d32297ab48da06934002068,
104'hb8659177cb2d3b395a00000000,
104'h90705591e0dc3c8eb8ac691f58,
104'h00fc52a8f8e7652ecee3b7d7c6,
104'h9c9b69583622f71d4502611804,
104'h54a63f864ce00e38c000000000,
104'h2c5c1c49b87a12a5f400000000,
104'h66565ebfacb64a166c00000000,
104'hbcd1c7f2a31460472800000000,
104'h94788fbbf1907e422000000000,
104'h305efc9dbd7f48dbfe00000000,
104'h0078f6a7f109ddf71382d49f04,
104'h3021cd5743d3a8fea700000000,
104'h28102871206da633db00000000,
104'hb86edbebddda6d0eb400000000,
104'h668016c4007c19aff800000000,
104'h345b24e7b6c0ed268100000000,
104'hbcadbc0a5bb53ce86a00000000,
104'hbc208b9541b909227200000000,
104'h54c3877287e5521cca00000000,
104'h28e92600d2a1049c4200000000,
104'h34c888e6916f1547deffffffff,
104'h084d48f99a8f22f41e00000000,
104'hbc585d15b08fb8221f00000000,
104'h9090540620dd0342ba4d57449a,
104'h9c67d967cf989e2a3100982201,
104'h30683d79d00ebc671d00000000,
104'h90c2780a84dad89eb518a09431,
104'h94dbde58b7b1b8f86300000000,
104'h90ac83e859c06276806ce19ed9,
104'h5483fe72070f53571e00000000,
104'h94d604b2ac4f1c719e00000000,
104'h543b2055764f319d9e00000000,
104'h288a6ace141189092300000000,
104'h90080d49106561a7ca6d6ceeda,
104'h34c8fb6c9121487b42ffffffff,
104'h90cf215a9ee8350ed02714544e,
104'h90b1fc7863cf54c29e7ea8bafd,
104'h901657592ca9dd3453bf8a6d7f,
104'h2874a09be925fd9d4b00000000,
104'hb8e814ccd0b1c7306300000000,
104'h94a9b3425340a4858100000000,
104'h04a0b60241f1b7e2e300000000,
104'h54c7049c8e3538b56a00000000,
104'h0832da0965d2a7e2a500000000,
104'h001795932f0b732d162308c045,
104'h942e6eab5c755f8fea00000000,
104'hb86483d1c9fdd2a4fb00000000,
104'h30967c702c42d3038500000000,
104'hb83ab5c37500579b0000000000,
104'h3451b2aba3283e1b5000000000,
104'h30794697f249004b9200000000,
104'h34c1b364839b007036ffffffff,
104'h3094b238295604b1ac00000000,
104'h04cd1f669a4039658000000000,
104'h08bac15075add2865b00000000,
104'h08686243d0d4240ea800000000,
104'h60c335508654c94da900000000,
104'h94693e3fd2ad334e5a00000000,
104'h0899345e32b4b63c6900000001,
104'h2831186b62f6edbced00000000,
104'h2889756a12721051e400000000,
104'h947a0491f48089b60100000000,
104'h66a12c1e426af447d500000000,
104'h9452913fa5bb49587600000000,
104'h9c09b4e913dbe09ab709a08813,
104'h941453bf2844967f8900000000,
104'h340d00f31a663189cc00000000,
104'h08e1341cc217dec32f00000001,
104'hb82ec2295d745d0de800000000,
104'h08f37926e6442f858800000001,
104'h288657380c37eee36f00000000,
104'h08cc946699c191dc8300000000,
104'h2c45778d8a3d44877a00000000,
104'h660eae2b1dc226aa8400000000,
104'h94179f512f510933a200000000,
104'h608cf17c199b02863600000000,
104'h00c63b728c3371e566f9ad57f2,
104'h94de9828bd20c9cf4100000000,
104'h084d959d9b55395baa00000001,
104'h0080b6bc01140c9f2894c35b29,
104'h604e803d9d9a5c0c3400000000,
104'h2c52c883a5f962d2f200000000,
104'hb888c27c11de9438bd00000000,
104'h66f9fb86f3794805f200000000,
104'h60ca444894b795da6f00000000,
104'h54773c97ee23b7954700000000,
104'h347efa4ffdb10aac6200000000,
104'h30fc033cf833889b6700000000,
104'h66cd91f89bfe4e2efc00000000,
104'h28c9ddc693ad89f65b00000000,
104'hbcecdd72d95de999bb00000000,
104'h9ca8bd3c51f75e40eea01c0040,
104'h541dffab3baacfea5500000000,
104'h6640017180c217d68400000000,
104'h3077584bee5759ddae00000000,
104'h285e44e9bce494d4c900000000,
104'h666c2fc1d8ce01ec9c00000000,
104'h54fbe8f4f7819b140300000000,
104'hbcbd23367a73e057e700000000,
104'h288461a00895b4362b00000000,
104'h603d50997ac8e7169100000000,
104'h00b241b664c8c994917b0b4af5,
104'h0898429430e1dde8c300000001,
104'h340a06c3141f80493f00000000,
104'h00049c9509381e47703cbadc79,
104'h00bfa5107fe85530d0a7fa414f,
104'h9c8f86c61f8b0f70168b064016,
104'h2c92d3ae250078eb0000000000,
104'hb86cda13d94f625f9e00000000,
104'h66ee1866dc4c6bcf9800000000,
104'h2c780c2bf0e80dd0d000000000,
104'hbc5493c7a90059fb0000000000,
104'hb8d1db74a3a50a3e4a00000000,
104'h08ea8d18d51437492800000001,
104'hbc46bb218d43cde78700000000,
104'h30a4be6849ff9b58ff00000000,
104'h04e9ff1ad36d88c5db00000000,
104'h346a6085d4995d843200000000,
104'h2811c80b236f2093de00000000,
104'h2835f6f76bb6f0e66d00000000,
104'h349faf603f26ecd14dffffffff,
104'h0400dc0d01e7805ccf00000000,
104'h9442334984e432b6c800000000,
104'h60058cd10b66ca85cd00000000,
104'h281ae2ad35b461446800000000,
104'h66a4b50e4923bdb74700000000,
104'h90f54938ea5a0d33b4af440b5e,
104'h28f8fb54f176d411ed00000000,
104'h90fa9b58f5e9acfed31337a626,
104'h60e58ceccbe42f6cc800000000,
104'h048e223a1cc814e49000000000,
104'h662b69e35605756b0a00000000,
104'h60be67ca7c86b2e00d00000000,
104'h94d17104a2776b65ee00000000,
104'h607722b1eed98aaeb300000000,
104'h54eb2bdcd6675275ce00000000,
104'h2c5fe25fbfa2f1c84500000000,
104'h288a5ab8141c03793800000000,
104'h9c137afb26d10b6ea2110a6a22,
104'h546740a1ce96cb0c2d00000000,
104'h081c3175388904981200000000,
104'h948baf661728058f5000000000,
104'h00e0a776c1dc1004b8bcb77b79,
104'hb80cd39119937b142600000000,
104'h666d876fdb0222310400000000,
104'h289fc06e3f207b814000000000,
104'h90c7f0868fd66d54ac119dd223,
104'h6094bc0c29b1ba6c6300000000,
104'h5434a2ab69119d6d2300000000,
104'h9c854b340ac0eb3481804b3400,
104'h609fea883f7dd439fb00000000,
104'h94c0fd7281da1cf2b400000000,
104'hbc124d8b242065334000000000,
104'hbc44f91389f2d684e500000000,
104'hbcddf5dcbb1551952a00000000,
104'hbcca472294b8f2867100000000,
104'h54f0de6ce198845e3100000000,
104'h9c36df6d6db53b546a341b4468,
104'h3477bee5ef78ce49f100000000,
104'h047d747ffaddc70abb00000000,
104'h04bdb7b27bf0a1d0e100000000,
104'h94b7ffa26ff41384e800000000,
104'h00f4be00e9a08f3241954d332a,
104'h00090ce512cae25e95d3ef43a7,
104'hbc52c7bba527806b4f00000000,
104'h2c8fc7121f4fd4f39f00000000,
104'h30afb78e5f94b5342900000000,
104'hb87ac3b7f5f4c860e900000000,
104'h049008e620af7f0a5e00000000,
104'h2c058f1f0bd4f180a900000000,
104'h30483bef90d0bd2ca100000000,
104'h30ecf854d9b1b8f06300000000,
104'h90a501944aca1892946f1906de,
104'h04a61d244ca3570c4600000000,
104'h084427838816fffb2d00000000,
104'h5464361dc8192ff13200000000,
104'h948a4426145363e1a600000000,
104'hbcb922867285ef780b00000000,
104'h54e122aac2b432806800000000,
104'h905cb46fb9d36540a68fd12f1f,
104'h34aaeefa55fd93d6fbffffffff,
104'hbc66bca3cd7a20a3f400000000,
104'h2c1621c52c32e59f6500000000,
104'h9007d6ad0fd8ccbeb1df1a13be,
104'h28be2c727cfc7754f800000000,
104'hb88cf4da19274c6d4e00000000,
104'h28c4e532897f0633fe00000000,
104'hbc39ac377321964b4300000000,
104'h90d0b2eca120f93741f04bdbe0,
104'h0445408d8a4650b58c00000000,
104'h661b795336795d1ff200000000,
104'h340670690c452dc78a00000000,
104'h547e44cbfc64a063c900000000,
104'h9c1a011934f9075cf218011830,
104'hb825b6854bfb0f40f600000000,
104'h34100aa92009bb131300000000,
104'h285b306bb6e50fb4ca00000000,
104'h34ec03e2d811c64323ffffffff,
104'hb88ec12a1d491d799200000000,
104'h08838e5207e3a20cc700000001,
104'h548dd02e1b4f860d9f00000000,
104'h9c880244104adf499508024010,
104'h089289a425f7e4aaef00000001,
104'h04c6bac68d650295ca00000000,
104'h2c980a7630bc5e4c7800000000,
104'h54ec21a2d86e204ddc00000000,
104'h601f4c513e3e9db17d00000000,
104'h04d57b66aa9d388c3a00000000,
104'h9c50d19fa1fa8f52f5508112a1,
104'h943d735d7a6c5331d800000000,
104'h2c27118f4ebadd6e7500000000,
104'h084f67939e685bd5d000000001,
104'h040da40d1b4b2c019600000000,
104'h006d74d1da64bdd3c9d232a5a3,
104'h66212dc142a414c44800000000,
104'h603542a76aaec04a5d00000000,
104'h94fc0c1af88ce3341900000000,
104'h088f8f601f9ca2143900000001,
104'hbcbbc146776f1091de00000000,
104'h90567c09ac9475ce28c209c784,
104'h04ab202e56d77fd0ae00000000,
104'hb8de986abd66bdd5cd00000000,
104'h04bd387e7ae179b4c200000000,
104'h546eaf15dd98c8423100000000,
104'h08c502a48a8768b40e00000000,
104'h66725151e4facaf4f500000000,
104'hbc15cbc92b95550e2a00000000,
104'h30f3232ae6a5bf864b00000000,
104'h04f861dcf0b920be7200000000,
104'h54a4e770493cff537900000000,
104'h0020ff8941ec837ed90d83081a,
104'h08904bac200f9f791f00000001,
104'h2811f8392334c6cf6900000000,
104'h2c28742d50758cd1eb00000000,
104'h901724192e7441e7e86365fec6,
104'h345747fbae8467f80800000000,
104'h34460c178cc995c69300000000,
104'h28cc7ce298f8214cf000000000,
104'h00aed5dc5db8a92671677f02ce,
104'h2c9b637236eb54e8d600000000,
104'h2ca9efd8531964853200000000,
104'h9cf372f4e6bb66a876b362a066,
104'h04ee7d34dc882e1c1000000000,
104'h047f9575ff345e296800000000,
104'h54dd81dcbbd425eaa800000000,
104'h66b833c070e082c2c100000000,
104'h082dce7f5ba721aa4e00000000,
104'h043401636817b7972f00000000,
104'h34e4ac84c96368d7c6ffffffff,
104'h30c388a6872a977d5500000000,
104'h90474a1b8ef330aee6b47ab568,
104'h08e3769ac6c551128a00000000,
104'h0430e62f6105d82b0b00000000,
104'h04d1a70aa36642b5cc00000000,
104'h04f9bc6af3f6e408ed00000000,
104'h3050f07fa184567e0800000000,
104'h2cdab13cb55abac7b500000000,
104'h2ce7b046cfc11e4c8200000000,
104'h9c79bdcff3ed209cda69208cd2,
104'h0825166f4a42afbb8500000001,
104'h2c0b1c0d165d7387ba00000000,
104'h943931bf721140232200000000,
104'h043332a56634a7456900000000,
104'hbcebbbc8d71480a52900000000,
104'h009541002ad10150a2664250cc,
104'h90bda4d27b0cba1919b11ecb62,
104'h34bacb4c753394e567ffffffff,
104'h34c15fec82a3a91c47ffffffff,
104'h66bfc6767f1b7f013600000000,
104'h6075eee1eb711a0de200000000,
104'h66ef842adfaae25c5500000000,
104'hbcb0ae3c618f45041e00000000,
104'hbc3e5ed17c91a3762300000000,
104'h5461e14bc31ae9e13500000000,
104'h284c25999879e48bf300000000,
104'h28bffe167fbb2c3a7600000000,
104'h305b486db63241956400000000,
104'h2825b96f4b0d2f731a00000000,
104'h6068c3fbd1d1cc50a300000000,
104'h54aed2dc5d8f72a01e00000000,
104'h0450cdada1d1c838a300000000,
104'h345fa0afbf68eca5d100000000,
104'h90ac3fb058d9268cb275193cea,
104'h94635befc627e8174f00000000,
104'h08d2c4eea5b5c2446b00000000,
104'hb8ad2c685a549f55a900000000,
104'hb82dc5195bbf5c1e7e00000000,
104'hbc07f4ab0f73987be700000000,
104'h08c8109490a056964000000000,
104'h9460ddffc1d3c164a700000000,
104'h28c64c928c4031e98000000000,
104'h54d8a470b1444bad8800000000,
104'h00341eff684bc811977fe710ff,
104'h04e7a2cecf8e48b21c00000000,
104'hb8521a81a49748ca2e00000000,
104'h28a09ea2414e058f9c00000000,
104'h34506a89a055f593ab00000000,
104'h94de5438bc8827201000000000,
104'h08223f4344e39da2c700000000,
104'h54e7c29ecf1686012d00000000,
104'h60d5f998ab9bd9fa3700000000,
104'h60d737a0aec8ca8c9100000000,
104'h289e17363cfb0952f600000000,
104'h9cd01bc6a0d4c8e0a9d008c0a0,
104'h9476de89ed050c290a00000000,
104'h60cf7e609ef29cd8e500000000,
104'h0414cabd29adc0b85b00000000,
104'h34a3617a4640860f81ffffffff,
104'h9c87b7be0fbf3efe7e8736be0e,
104'h9454c5dda9ca83e29500000000,
104'h54bece367d79d4b5f300000000,
104'h2c1077192051b16da300000000,
104'h54d92f96b2e9c15ad300000000,
104'h305a9775b5af618c5e00000000,
104'h34ef6204deaeb22a5dffffffff,
104'h9c18ec0131effadadf08e80011,
104'h30c17c7082b0fe1e6100000000,
104'h04bfe8867f0193b50300000000,
104'h54761285ec00a1f50100000000,
104'h60ae7b945c924e362400000000,
104'h3055e0afabd9fc28b300000000,
104'h34849a74097a743df4ffffffff,
104'h94303819608c48f61800000000,
104'h30008d3301ce53609c00000000,
104'h66d42aaea8bdde5a7b00000000,
104'hbcaefa9c5d73d903e700000000,
104'h00ca771e944a281194149f3028,
104'hbc79b43df3d7ee3aaf00000000,
104'h903c34d378b563946a89574712,
104'h54e14260c21f93e93f00000000,
104'h00b23ff664f21c20e4a45c1748,
104'h006d3013daf0bea4e15deeb8bb,
104'hbc19657932f466b2e800000000,
104'h549f171e3eaef2cc5d00000000,
104'h66374f036e4ede099d00000000,
104'h9c746c13e8c7a07c8f44201088,
104'hbc7c2f03f8d55e9aaa00000000,
104'h00430a39866a3f91d4ad49cb5a,
104'h34dd2ca2ba0182a703ffffffff,
104'h347c7f9df8c82ba29000000000,
104'h60238fcf4794de282900000000,
104'h90a4190c48b84012701c591e38,
104'h28dcad34b9b4fada6900000000,
104'h0483ae12075a33f9b400000000,
104'h9cd6923ead7d143dfa54103ca8,
104'h9c6b2cfdd615b6352b01243502,
104'h34d57118aac1938683ffffffff,
104'hb806e6d30d11495f2200000000,
104'h54edccb0db814bb80200000000,
104'h2c189b6731fcdfd4f900000000,
104'hbcaf64b05e40758b8000000000,
104'h901f453f3ecc37b298d3728da6,
104'h900ce18719496b7b92458afc8b,
104'h00b9a5aa73bcf6d279769c7cec,
104'h66ac405c588f25c41e00000000,
104'h9c4f90b79fc486d48944809489,
104'h300bff1f17ad76645a00000000,
104'h2c4df92d9b41b1138300000000,
104'h34a9087a5243051786ffffffff,
104'h5401bc99038dfaa61b00000000,
104'h2c115fdb22a10b544200000000,
104'h08dd2f46bacac06e9500000000,
104'h908f8d6c1f8cd05e19035d3206,
104'h66b46844680613090c00000000,
104'h54daca18b58ee52c1d00000000,
104'h083c4d5d789352cc2600000000,
104'h60f7eb90ef0c207f1800000000,
104'h04d85f1cb0338bd96700000000,
104'h3037103b6e245acd4800000000,
104'h9c8344ce06699207d301000602,
104'h60fa0b46f412ea552500000000,
104'h085e187fbc15dcf72b00000000,
104'h54af90a05f8cdf121900000000,
104'hbc3272fb643624036c00000000,
104'h082f20f15e58fec1b100000001,
104'h30f337cce664ba45c900000000,
104'h9061b5a7c31d80df3b7c3578f8,
104'h540821431073aa9be700000000,
104'h28e32ceec61f8aa53f00000000,
104'h34f00c66e03f93a37fffffffff,
104'h000875b310706b13e078e0c6f0,
104'h2c8605040c9643b42c00000000,
104'h9c767b9fecc496e08944128088,
104'h94f511aaeacd14ee9a00000000,
104'h2835d31f6bf0648ce000000000,
104'h0826bfa34d63092bc600000001,
104'h90ef2560dec688528d29ad3253,
104'h9c386ef970caa6089508260810,
104'h04bc5c5078d4502ea800000000,
104'hbc435e7b863790e36f00000000,
104'h94ba8e9675379fdd6f00000000,
104'h288377b2060bead31700000000,
104'h0048aba5918aacd615d3587ba6,
104'h28a8daee51416cb78200000000,
104'h049ee7a03da17a5c4200000000,
104'h66e02b36c0ea432ad400000000,
104'h002ae77b559515662abffce17f,
104'h60dd9a5cbba5aa8c4b00000000,
104'h08dcacdcb95890b3b100000001,
104'h54f6b4e6eda44af24800000000,
104'hb8504235a0d3c0bea700000000,
104'h6016ee252d98543e3000000000,
104'hbc8026ac003fb7c37f00000000,
104'hbc1aec2335ad5a0a5a00000000,
104'h286c7a31d84101bb8200000000,
104'hb8de93aabd63efb3c700000000,
104'h34e2e96ec5fba066f7ffffffff,
104'h9009d44913ed0450dae4d019c9,
104'h005359d1a61cc74139702112df,
104'h66683449d060fec3c100000000,
104'h605d5583ba9657822c00000000,
104'h94571cb9aeee99a4dd00000000,
104'h9482377204881c2c1000000000,
104'h2c96e5622ddd7f52ba00000000,
104'h3028174b5092c5f62500000000,
104'h048aa0d41500a5e90100000000,
104'h28d97578b290a75e2100000000,
104'h34b2a85865f46b42e8ffffffff,
104'h546da727db7030a1e000000000,
104'h2cede7fadb4470fd8800000000,
104'h908602400cac2bb8582a29f854,
104'h54cdea889b553871aa00000000,
104'hb88bc974179db8623b00000000,
104'h5409a58d13ad7ebe5a00000000,
104'h901ad82d35a4081848bed0357d,
104'h94db0554b6fb58bef600000000,
104'h9c850e940addda1abb850a100a,
104'h28d338eaa6f10f0ee200000000,
104'hbcda7d9ab4f0b760e100000000,
104'h3071be1be3d5ba0aab00000000,
104'h60a252e84419eea93300000000,
104'h048a2d7214659dcfcb00000000,
104'h003084ed6185506e0ab5d55b6b,
104'h0044c63d895e4637bca30c7545,
104'h34443ed188a5aaee4b00000000,
104'h9045ba858bd262dea497d85b2f,
104'hb85b0c81b60b06251600000000,
104'h9c473b198e2163214201230102,
104'h94e4c6aac9f29fcce500000000,
104'h28324383642ed21d5d00000000,
104'h08443eb9888ca7621900000000,
104'hbc822610043572ab6a00000000,
104'h3048aad991b3ba206700000000,
104'h007ed7cdfd521b69a4d0f337a1,
104'h9c8bd1f217921f042482110004,
104'h5499fc8233a252b24400000000,
104'h60e0f7b8c170c2cde100000000,
104'h94fab2bef592aaa42500000000,
104'h94c0889081abf3f05700000000,
104'h04041fcf08b8dd1a7100000000,
104'h665c85abb989deae1300000000,
104'h3462bbbfc555a7b1ab00000000,
104'h2cc9b0f0936ec903dd00000000,
104'h90ec5d58d85a67c1b4b63a996c,
104'h9c697911d2ab0ea65629080052,
104'h905f0629be8e766a1cd17043a2,
104'h0880a57401dedd1abd00000001,
104'h00ca6e7a9430448760fab301f4,
104'h28a6c24a4dafaf985f00000000,
104'hb830515d602e36b35c00000000,
104'h907a4c7df44b8b1b9731c76663,
104'h08a778984ed3414aa600000001,
104'hb8c59db68bf5fa5eeb00000000,
104'h280d88bd1b83446a0600000000,
104'h94009865019ac9e03500000000,
104'h60138d1327e327eec600000000,
104'h2cdb13b4b62283dd4500000000,
104'h343143a96288b7721100000000,
104'h303c07937804ac4f0900000000,
104'hbccb2946960e3e511c00000000,
104'h66e178a6c253bcf3a700000000,
104'h5497457c2e25e3a94b00000000,
104'h668d24601a3ee1437d00000000,
104'h940cb6971908c6531100000000,
104'h2c69ecedd3c5727e8a00000000,
104'h9469fd9fd35dd8edbb00000000,
104'h901605352c18339f300e36aa1c,
104'h2c9e0a603c747dd3e800000000,
104'h047ddce5fbe44d62c800000000,
104'h9c20076b406ee321dd20032140,
104'h9473cc6be7840a420800000000,
104'h3481e60603b81eb270ffffffff,
104'h04b080ee61d1527ca200000000,
104'h6049aa4193e20a24c400000000,
104'h04a828625015e80d2b00000000,
104'h305d76e7bac6ded08d00000000,
104'h04605d6fc05562adaa00000000,
104'h600e59831c8a91d61500000000,
104'hb832d37f65ecebdcd900000000,
104'h9c8dd6621bd7f00eaf85d0020b,
104'h2c28c2bf5144bad58900000000,
104'h545a3491b4757a17ea00000000,
104'h305b141db60f50951e00000000,
104'h54ed89d8db0e004b1c00000000,
104'h30834d42065273d5a400000000,
104'h34bb86c877c8fec691ffffffff,
104'h28a93c9e5235ed136b00000000,
104'h664a02ab940eb9671d00000000,
104'hb899655a3254028ba800000000,
104'h9cf0478ae09417c62890078220,
104'h94902b622007b4390f00000000,
104'hbc891e36128a41401400000000,
104'h2c45bf658bf4b7d8e900000000,
104'h2c239a39478df8f41b00000000,
104'hb846cacb8dc534e48a00000000,
104'h087ea5ddfdb2b9ba6500000000,
104'h3045dbc18bd9409cb200000000,
104'hb8db4e30b6c592308b00000000,
104'h00d19134a36419f9c835ab2e6b,
104'h9471cf01e3a3c0b24700000000,
104'h669b86d0373325b76600000000,
104'h9c955ed42a410f5d82010e5402,
104'h083c0103781aaa553500000000,
104'h2852bafda5b9f00a7300000000,
104'hbc1e58f53cc44c0a8800000000,
104'h2c1573852a8d58581a00000000,
104'h08022893045b48d5b600000001,
104'hbc9ff7343fda5da0b400000000,
104'h283d368b7a527473a400000000,
104'h00625f9fc43d91037b9ff0a33f,
104'h34aa2246543ff45f7fffffffff,
104'h08fbfd08f7aa1b565400000000,
104'h66efcff2df8abbd21500000000,
104'h5473a283e75a993bb500000000,
104'h668d947c1b65c7cfcb00000000,
104'h0072b1d7e5b5b70a6b2868e250,
104'h90d82190b0551b0baa8d3a9b1a,
104'h2c8ee7921dc28ce28500000000,
104'h60d33196a6387a057000000000,
104'h906ee701dd88ba9e11e65d9fcc,
104'h2c93f3be2797e6f82f00000000,
104'h2855862dab7843d9f000000000,
104'h9c9837f230addde25b8815e210,
104'hbc5fd9e5bfb52bf06a00000000,
104'hbc3e5ae17c6b507fd600000000,
104'hbc8201b204e2d1fec500000000,
104'h0849f1f393716247e200000001,
104'h900eb3e51dcb0ce296c5bf078b,
104'hbc21375742bce47a7900000000,
104'hbc558985abfd0734fa00000000,
104'h082f35f55e7f9213ff00000001,
104'h60a40a5e483fdb537f00000000,
104'hb896b57e2d630bcdc600000000,
104'h04b579006a74ef59e900000000,
104'hbc21e65b433194256300000000,
104'h045d5eb5ba4611238c00000000,
104'h661acdb935a08b564100000000,
104'h54f8d786f1bb524a7600000000,
104'h94787185f0b8ab5e7100000000,
104'h94f29e44e594a4302900000000,
104'h9c8cc466191803f93008006010,
104'h6665d879cb0333ed0600000000,
104'h901f51cf3e09b6a11316e76e2d,
104'h66aba26e571e865f3d00000000,
104'h2ca0a9e8412f72915e00000000,
104'h2c5f5b35be31541f6200000000,
104'hbce28d9ec538b0c97100000000,
104'hbc25b0974bba258a7400000000,
104'h0880da9c01e3b000c700000001,
104'h2c426b1d84bbaebe7700000000,
104'h9ce7374ece4430b78844300688,
104'h54c8fa1691b8eb967100000000,
104'h049f7ee23e0bf1271700000000,
104'h54f3bf90e778fbadf100000000,
104'h0854ed45a950e94da100000000,
104'h30ee1c52dc6ebe61dd00000000,
104'h04b80b1c700d46e31a00000000,
104'h541d3bef3a602ecbc000000000,
104'h002f59dd5e552969aa84834708,
104'hbcb3a0aa67a97fca5200000000,
104'h0400bfab01fe1e18fc00000000,
104'h541b6f973637f7f96f00000000,
104'h665fb377bf345bed6800000000,
104'h60837c7c06188db33100000000,
104'h9c8c28ea1839bfa3730828a210,
104'h089b15ea363643156c00000001,
104'h66ee3c74dc4a87b79500000000,
104'h6648912b91a441fa4800000000,
104'h04da9f3eb563d065c700000000,
104'h04e69648cd8fb7fe1f00000000,
104'h346bc335d767cfa9cf00000000,
104'h90542c13a8b572806ae15e93c2,
104'h949bc70437dbd13eb700000000,
104'h04e38412c7f73a98ee00000000,
104'h9c8b2218163bf2a3770b220016,
104'h54f38696e76cf127d900000000,
104'hbca0109c40a09f0e4100000000,
104'h54c01ea8800d6ac31a00000000,
104'h9ceabf7ed531cb8163208b0041,
104'hb8b546146acb0bca9600000000,
104'hb8fa3868f4a3f2b64700000000,
104'h6650d169a1c0245a8000000000,
104'h600e0dc91cbad1287500000000,
104'h045efbefbdc70c4e8e00000000,
104'h6050c6c9a18de1141b00000000,
104'h9c1db3b33b99ff403319b30033,
104'h2c870b540e0a96771500000000,
104'h6092a5822556b891ad00000000,
104'hbc5f901bbff05b08e000000000,
104'h9c2008e94001cf570300084100,
104'hbc4fc2859f424a4b8400000000,
104'h04242c334865d273cb00000000,
104'h60a934be52eaad74d500000000,
104'h042fc0695f6a247dd400000000,
104'h0453c9b7a70c37871800000000,
104'h2c1ee55d3dbd97d27b00000000,
104'h9058a117b13d01397a65a02ecb,
104'h0020f5954170ca91e191c02722,
104'hbc29c34d53a745084e00000000,
104'hbc7b1261f6dc4290b800000000,
104'h66528d83a5cbdb329700000000,
104'h08916fcc22ee4972dc00000001,
104'h9cfcdda4f96275b3c46055a0c0,
104'hbc8360a206bc88907900000000,
104'h9c76fe61ed939c4427129c4025,
104'h2c66226fccf56504ea00000000,
104'h04a653204c8868621000000000,
104'h60ea697cd48d1bac1a00000000,
104'h6612c413250c014d1800000000,
104'h34f8acdaf1c29d2685ffffffff,
104'h34f6ea1eedbad7fa75ffffffff,
104'h00903252205829cbb0e85c1dd0,
104'h5480faf601fba32cf700000000,
104'h66f4da72e99badb63700000000,
104'h0430750160be1b5a7c00000000,
104'h28f7ac84ef9adcc43500000000,
104'h66fc8b6cf9bb76c27600000000,
104'h08e62294cc9f0e943e00000000,
104'h94af52265eb4a5606900000000,
104'h006c3571d8ccda8099390ff271,
104'h00a1a9d643ea4ceed48bf6c517,
104'h287528a3ea8373a20600000000,
104'hb8c3ebec87ca84ec9500000000,
104'h2cd71678aed7c4d8af00000000,
104'h089f56943e9052922000000000,
104'h04553bfdaa474cc18e00000000,
104'h9cbc38b87850e4e1a11020a020,
104'h604504fb8a7eb9b3fd00000000,
104'h0098de0431b2908e654b6e9296,
104'h54e1d800c3d045cca000000000,
104'h301d3ae53a498c1b9300000000,
104'hbc1ba25937b5d2e86b00000000,
104'h603758876e566bc1ac00000000,
104'h546c240fd87ac6a7f500000000,
104'h600c80d719625d7dc400000000,
104'h94fefbf0fde9a660d300000000,
104'h94eb2a7cd6f5250aea00000000,
104'h66387389709973303200000000,
104'hbce9a4ead360d7e5c100000000,
104'h94670b25ce36c5f56d00000000,
104'h54dd8446bb5f594bbe00000000,
104'h082bc5cd57e4ab48c900000000,
104'h0817cd812ffd9634fb00000000,
104'h2ce53552ca913f8a2200000000,
104'h2c11e243231081612100000000,
104'h0029463d52da0ad0b403510e06,
104'h30f72cfaee2fcf4d5f00000000,
104'h6019cbdb33dc1cfcb800000000,
104'h9cb78cd26ff27230e4b2001064,
104'h281fcc393f0be9a91700000000,
104'h340e81b71de8d608d100000000,
104'h60598c21b3f0e430e100000000,
104'h28ab18545690dc942100000000,
104'h66c75b1e8e60dbafc100000000,
104'h30649617c93f994f7f00000000,
104'hb8031f7f069717002e00000000,
104'hb827e5294fbccd707900000000,
104'h9c0ea24f1d4330c38602204304,
104'h9409c079130c23fb1800000000,
104'h00849b58096bb351d7f04ea9e0,
104'h9ca99fb053a02da440a00da040,
104'h04387d2b70c074c68000000000,
104'h00d1633ea2f31cece6c4802b88,
104'h5411010f22b8b3007100000000,
104'h04fdc04cfb41420f8200000000,
104'h54a973105298ef9a3100000000,
104'hb83b6cc776e14706c200000000,
104'h3005bdff0b3c8bef7900000000,
104'h94850b5a0a762b91ec00000000,
104'h34653763ca3f251d7e00000000,
104'h908dd7721bf70126ee7ad654f5,
104'h30002b8b00e1affcc300000000,
104'h08a5113a4a4867099000000001,
104'h343c298178c7552c8e00000000,
104'h041e29a13ce3c62ec700000000,
104'h60a30f1046660d09cc00000000,
104'h3469ae4fd3c84d569000000000,
104'h94a8d4c851c6fbac8d00000000,
104'h2ccaf5b295b1acfc6300000000,
104'h340c19f318f28cf4e500000000,
104'h66568af7ad50935da100000000,
104'h305d709bba24507d4800000000,
104'hb8a55a064a00e8730100000000,
104'h00f9698ef2a2959e459bff2d37,
104'h04689b91d139c9fb7300000000,
104'h9c81605802d5c77aab81405802,
104'h30ca80fe95b347706600000000,
104'h089f07463efb88e8f700000001,
104'h9047a07f8ffdde0efbba7e7174,
104'h349eb3623d91908623ffffffff,
104'h286d20f9da07b4d30f00000000,
104'h002c6879585444b1a880ad2b00,
104'hb8a7a61e4fcb987a9700000000,
104'h543fa5157f6d1783da00000000,
104'h080efc571d25b77f4b00000001,
104'h9c01ee85032ca2d95900a28101,
104'h9cda84d0b58a1e1c148a041014,
104'h083c1cd5786c844fd900000001,
104'h66ea6176d418f2513100000000,
104'h2c9666ce2c74f93fe900000000,
104'h089160f6224c6fd59800000001,
104'h30b72dfe6e023ac90400000000,
104'h288baaba173ca4297900000000,
104'hb80c8ab119c599c48b00000000,
104'h94ce2af09c34ea876900000000,
104'h66cc97f2997e5ad1fc00000000,
104'h549abe82351727e92e00000000,
104'hb8787f8ff08652480c00000000,
104'h34051f1d0ac8c70c9100000000,
104'h60ee4612dc6e4049dc00000000,
104'h28d48f2aa9a5746e4a00000000,
104'h08d556c8aa05ecad0b00000001,
104'h086e45dbdcb39a4a6700000000,
104'h28f1cfbee3ec0310d800000000,
104'h08349b1969169c9d2d00000000,
104'hbcaa8dbc5581aece0300000000,
104'h6686f38c0dfad520f500000000,
104'h94cdf8529bddf706bb00000000,
104'h944e6ca79cf74f50ee00000000,
104'hbc618dcdc31cda913900000000,
104'h2cc3489286a1446c4200000000,
104'hbc082f3510262c0b4c00000000,
104'h9cd71a3aaecd576c9ac512288a,
104'hb84b2c5796c82dd09000000000,
104'h2c6fb14bdfba91107500000000,
104'h60d20fc0a4c1edfe8300000000,
104'h285ec631bd231bd14600000000,
104'h66552abdaa1962713200000000,
104'h00c2661484eebfeaddb125ff61,
104'hb8d6e156add944c2b200000000,
104'h283a1ee974031f5b0600000000,
104'h046fb65ddf12ae4f2500000000,
104'h081ceb55396db1dbdb00000001,
104'h90b9175872be74347c07636c0e,
104'hbc9bdec437e380eac700000000,
104'h08a2e89845da434cb400000001,
104'h2c7d9165fb52a3c3a500000000,
104'hb83fd1277fdd7c34ba00000000,
104'hb8de4c22bc017b630200000000,
104'h60d446cea861cf49c300000000,
104'h3020f4a94177ae83ef00000000,
104'hbc345a1f689b98a43700000000,
104'h94fcb964f92ce5a15900000000,
104'h663c426178fdfc24fb00000000,
104'h94537d81a6b946f87200000000,
104'h54efa9a0df26c1654d00000000,
104'h603d04e97a03b2870700000000,
104'h008bb8ac17edefbedb79a86af2,
104'h6072e04be5a9be065300000000,
104'h9097e30e2f352a536aa2c95d45,
104'h9c091911129d70f23a09101012,
104'h34c1731282d2cbf8a5ffffffff,
104'h541f9d673fb4c08a6900000000,
104'h300dd5c71bb4c34e6900000000,
104'h00f86c3af0a6cbc64d9f38013d,
104'h66afa6f65f172eb12e00000000,
104'hb89e81363db2d7646500000000,
104'h2c8a7d2a146ab83bd500000000,
104'h000980c913ed09e2daf68aabed,
104'h343175b36246b1c98d00000000,
104'h906a241bd4ece778d986c3630d,
104'hbcec809ad982f0f60500000000,
104'h600b651916598e23b300000000,
104'h04106cab20556b1faa00000000,
104'h60f46a70e88fb1a01f00000000,
104'h08b5b3746b0f91611f00000001,
104'hb837338d6e5d576dba00000000,
104'h289a053e34d76c94ae00000000,
104'h34980498308f52c01effffffff,
104'h34b8951871787959f0ffffffff,
104'h2cf99282f3cc809c9900000000,
104'h30e524ccca2844095000000000,
104'h90b9eef673fac3b8f5432d4e86,
104'h2875d0e9ebdac4c0b500000000,
104'h94ec345cd829c0935300000000,
104'h28c79cb68f827b5c0400000000,
104'hb81af1e535bf59667e00000000,
104'hbc29be4353584b77b000000000,
104'h9cff5778fe61ea31c3614230c2,
104'h307baa5bf707186f0e00000000,
104'h945921c7b2dc44acb800000000,
104'h2889e0881357215dae00000000,
104'h08d34638a6f76c54ee00000001,
104'h94f5771aeab51d206a00000000,
104'h00a15efc420612690ca771654e,
104'h0032671b64b1165262e37d6dc6,
104'h2841d6fb839dd1e03b00000000,
104'h30e89854d1510751a200000000,
104'h6690d5e421ba2b7a7400000000,
104'h00c3ad5687d33636a696e38d2d,
104'h2817ec212f4541b38a00000000,
104'h347d8f6bfb3c50e17800000000,
104'hbc467edf8cc254c48400000000,
104'h08afba9c5fcd48e89a00000001,
104'h28fef40afd95feac2b00000000,
104'h66b749ba6e3cefaf7900000000,
104'h08a49e4c49282f275000000001,
104'h2cb7c24e6f51524ba200000000,
104'h2c9669142cdbe7aeb700000000,
104'h6688a0a41134d59d6900000000,
104'h94c2448e8498b77e3100000000,
104'h0419a3cb33a3123c4600000000,
104'h30bd51a47a61f797c300000000,
104'h9c99d98c33c970889289508812,
104'h668cce021937c6af6f00000000,
104'h946d6a73da77849def00000000,
104'h540bc015173dc5457b00000000,
104'hbcbe25cc7cfb2a54f600000000,
104'h9099630832e39194c77af29cf5,
104'h0032cda765c4614a88f72ef1ed,
104'h667c52cbf88b039a1600000000,
104'h901922c932ace8de59b5ca176b,
104'h282678034ce82910d000000000,
104'h900eb0c51d7f9c29ff712cece2,
104'h9445b4238b1701772e00000000,
104'h90f459e0e81b8e0937efd7e9df,
104'h944d4d519a22fa074500000000,
104'h9cb8a32c714ee5179d08a10411,
104'h54e41a7cc87c29bbf800000000,
104'h5444c073894577b18a00000000,
104'h9c636f51c6964d502c024d5004,
104'h30986040302727f34e00000000,
104'h3452c83ba5ad83445b00000000,
104'hbce037e0c041ffb98300000000,
104'h548c3664186cc7d3d900000000,
104'h94134f5f26dc0c9cb800000000,
104'h54758bbbebf230f6e400000000,
104'h28630d89c688fbfe1100000000,
104'h947a46ebf46cea6dd900000000,
104'h348a03e8149f76f63effffffff,
104'h2cb23f5e6450f1b1a100000000,
104'h00c57acc8a2a3e6554efb931de,
104'h04611143c2dc91fcb900000000,
104'h9c05bd3f0b7106e1e201042102,
104'h94ba4984746ba04fd700000000,
104'h34a1250a42f514c8eaffffffff,
104'h301651cf2cd47764a800000000,
104'h9495e6be2b7d9839fb00000000,
104'h60841c8e08cab3b69500000000,
104'h9c269da54d8fc90c1f0689040d,
104'h9c6390efc703af830703808307,
104'h605d97c9bb6ec2dfdd00000000,
104'h2c74b6dbe998bec43100000000,
104'h90c2e1f8857f210ffebdc0f77b,
104'h3087a3000fe32b36c600000000,
104'h945113bfa2aa5ab45400000000,
104'h08b922ca72cdf0589b00000001,
104'h6674db69e91ddeb13b00000000,
104'h08e82864d0593763b200000001,
104'h30a349fe4681ef9a0300000000,
104'h2ccff6bc9fcb93549700000000,
104'h28d2df52a5843fd00800000000,
104'hbcf30d7ce6ccfce69900000000,
104'h34e355eac6524d6fa4ffffffff,
104'h5442d51385678e97cf00000000,
104'h94c02f16805f7e4fbe00000000,
104'h60300aa960aa00a05400000000,
104'h94c9fee29392fc102500000000,
104'h948fec2a1f67e501cf00000000,
104'h90d27818a4b9500e726b2816d6,
104'h008224460453a373a7d5c7b9ab,
104'h66b738446ed5bf62ab00000000,
104'h90437667866e3571dc2d43165a,
104'h9c6753b3ceaf66ea5e2742a24e,
104'h00992ab83288a23a1121ccf243,
104'h60dfa170bfb617446c00000000,
104'hb8413a2582533ac9a600000000,
104'h2869c749d31af0c93500000000,
104'h94933a5c263695db6d00000000,
104'h542a05c954b8bf947100000000,
104'h9c3e09c77cf24be8e43209c064,
104'h34c7c43a8f28178350ffffffff,
104'h9cce3b929cbd73307a8c331018,
104'h54bcdcaa791b30333600000000,
104'h2c6943add264dbafc900000000,
104'h2c97a7e62fdd80febb00000000,
104'h28e962bcd2a30b1c4600000000,
104'h083bc97977931d002600000000,
104'h304652338cadf8fa5b00000000,
104'hbcedbbaedb93cf162700000000,
104'h30f6b03aedb68a806d00000000,
104'h08b51b926afdf5defb00000001,
104'h00b62bbe6cd5ceaeab8bfa6d17,
104'hb861b4f1c35d1fb1ba00000000,
104'h2cdc706ab8a3fa3c4700000000,
104'hb83f4e577e0066ab0000000000,
104'hb830d2ab617523a9ea00000000,
104'h2c44350f885c8ca7b900000000,
104'h04e6bbaccdf7bf2eef00000000,
104'h084689258d95d7442b00000000,
104'h602ed55d5db0daca6100000000,
104'h30844966080dabdf1b00000000,
104'h0888f66211921a382400000001,
104'hbc8a1f5e148feb8e1f00000000,
104'hbcc2ce3085a572f24a00000000,
104'h9044eb5b897c0f33f838e46871,
104'h004f50ed9e8aa83815d9f925b3,
104'h9cca1062940603670c02006204,
104'h0862e387c54287038500000000,
104'h04228049456ac489d500000000,
104'h340047a90083e20e0700000000,
104'h3024879349b4baae6900000000,
104'h00e247c0c4964dda2c78959af0,
104'h54285991506bd5bbd700000000,
104'h2cee22f8dc6e9c9fdd00000000,
104'h04235c4f464d69479a00000000,
104'h9c9ab93c35891a561288181410,
104'h90763497ece7c8aecf91fc3923,
104'h0478773bf0bd88c27b00000000,
104'h607991f5f3b5a30c6b00000000,
104'h60c6025c8c08db5d1100000000,
104'h3095bab42b151f3f2a00000000,
104'h66bda4ce7b08b35f1100000000,
104'h9c70d7e5e136b7e16d3097e161,
104'h2807797f0ea49bc84900000000,
104'h9480014e00dfd74ebf00000000,
104'hb87c5817f82105534200000000,
104'h660709810e9d33a43a00000000,
104'h342581054b98027a3000000000,
104'h2c5309c5a6c0eabe8100000000,
104'h082509734a93c37c2700000000,
104'h54bbae2677485e399000000000,
104'h00f3074ce646d2558d39d9a273,
104'h04b741746e85cf6c0b00000000,
104'h941b7d41369e0ebe3c00000000,
104'h000d79391a29bb7b533734b46d,
104'h606906b9d2286a355000000000,
104'h94f501c0ea07f73b0f00000000,
104'h662843e1509063f62000000000,
104'h00a7ca164fb48b4a695c5560b8,
104'h2cf005a6e02344fd4600000000,
104'h2cba100674d45006a800000000,
104'h541a39b534a21c044400000000,
104'h66402c1f80bd498a7a00000000,
104'h00d99678b358798bb032100463,
104'h308f1da81ec2c3b28500000000,
104'h6698071c3034ebcb6900000000,
104'hb823d6b147492e1b9200000000,
104'hb809d78d135f3ac1be00000000,
104'h54fd4804fa7db81dfb00000000,
104'h0421a077438864281000000000,
104'h9c752d2fea4dacd99b452c098a,
104'h2cd0f344a1f0577ee000000000,
104'h9c63987dc7f98f26f3618824c3,
104'h0841c62583dd71fcba00000000,
104'h34193ef9325ff5a5bf00000000,
104'h08f49ffee901baa10300000001,
104'h667c846ff9dc26aeb800000000,
104'h00ef8484df09de2913f962adf2,
104'h9455476baa547461a800000000,
104'h00e9a01cd351eb0da33b8b2a76,
104'hb8936d3a26d45896a800000000,
104'h661fb3f73f7bcd8bf700000000,
104'h001c2deb38ce50ec9cea7ed7d4,
104'h303d41fd7a638b9fc700000000,
104'hbc6a2045d4e17abcc200000000,
104'h288678dc0cad41025a00000000,
104'h000c05d518beef267dcaf4fb95,
104'h082ee0015de8db36d100000000,
104'hbcce56e69c8adf021500000000,
104'hbc88c396110795750f00000000,
104'h2c1b8e8937d56eeeaa00000000,
104'hb8796089f29f34b63e00000000,
104'h28df3684be0753470e00000000,
104'hbc5dd083bb3703bb6e00000000,
104'h28f7b368efde2c26bc00000000,
104'h044cb5f1999a8efc3500000000,
104'h9002d07f0554a16ba9567114ac,
104'h9460a801c1ee20b8dc00000000,
104'h00110bd522123eaf24234a8446,
104'h54775e9fee00fceb0100000000,
104'h308ba232173f0f4d7e00000000,
104'h9c919e7223195d4f32111c4222,
104'h54595b29b256fa65ad00000000,
104'h00bfe4ec7f362d5f6cf6124beb,
104'h540e15031c58decfb100000000,
104'hbc47d4398f82865a0500000000,
104'h30b110ca626d6f29da00000000,
104'h906e5f41dc76eb3bed18b47a31,
104'h3065fe4dcbe1cdcec300000000,
104'h2c12b5b125e444bec800000000,
104'h0004c8170911e8dd2316b0f42c,
104'h6005eff70be49d5ec900000000,
104'h286c1f73d89e962e3d00000000,
104'h2ccb7b3a966d9d59db00000000,
104'h041ac86d350b6f611600000000,
104'h2c2e456f5c00c6a90100000000,
104'h345ba5d3b7a06dcc4000000000,
104'h2cd6a93aadb571086a00000000,
104'h2810852f212b46935600000000,
104'h94cd1a0a9a9885f83100000000,
104'h9ce7aacecffc868af9e4828ac9,
104'h9c95900a2b1dfcb13b1590002b,
104'h2c881dbc103c6e537800000000,
104'h944fb4299f2016314000000000,
104'h0000b3c501738e47e774420ce8,
104'h2807cc0f0fa859305000000000,
104'h9085dd740be32282c666fff6cd,
104'h2c24662b487e4e2ffc00000000,
104'h664a321794092ee31200000000,
104'h669cc5a63937fb676f00000000,
104'h28fdbbb6fb6c5b03d800000000,
104'h2c640e6fc84820d59000000000,
104'h90400323808b8e3c17cb8d1f97,
104'h903531316a4634358c730504e6,
104'h3410dbe5218d4bb01a00000000,
104'h60ab9756576c1d01d800000000,
104'h040bf049170ace371500000000,
104'h60548f0da905b0790b00000000,
104'h30fb0d5cf612e46d2500000000,
104'h002577414a4ded959b7364d6e5,
104'hb80b2eed16408caf8100000000,
104'h5482ab9c05f5f912eb00000000,
104'h04b04b80608151180200000000,
104'h34c3308e8651d971a3ffffffff,
104'hbc03e06907e76386ce00000000,
104'h54dd1f40bae6f2e6cd00000000,
104'h042a3db154a379944600000000,
104'h2ca6d19e4dd84370b000000000,
104'h300a92211502689d0400000000,
104'h34d8ce56b16c5ecfd8ffffffff,
104'h9465b74bcb0a81bf1500000000,
104'h34bc74d278a92a7a52ffffffff,
104'h0817bd752f14add32900000000,
104'h2833693f66c159ae8200000000,
104'h901037af207d4977fa6d7ed8da,
104'h6683c08807cfa96a9f00000000,
104'h9c4d47c39a48c1079148410390,
104'h0814ec5d291bdc673700000001,
104'h04e56a3eca57ec9faf00000000,
104'h3009672312e57720ca00000000,
104'h00ec026cd8882c1a10742e86e8,
104'h9061200bc2703bd5e0111bde22,
104'h54bca65879db4314b600000000,
104'h9410a6ff21ce667e9c00000000,
104'h30f92ad0f282f4ec0500000000,
104'h543918ad72a4a8da4900000000,
104'h2c466f5f8c6c60bbd800000000,
104'hb86cca7fd9e3e662c700000000,
104'h9093ea5027a71d5e4e34f70e69,
104'h34acb6a25934b05769ffffffff,
104'hb879f4b1f3c415708800000000,
104'h2c8aa800159081ae2100000000,
104'h66fad64af508234f1000000000,
104'h909c264a3844bb2989d89d63b1,
104'h28b291ac650e6d151c00000000,
104'h902a21e7545b5f41b6717ea6e2,
104'h344170218236809f6d00000000,
104'h34c9600492258e334bffffffff,
104'hb87d4db3fafa2f86f400000000,
104'h3047a6918f63c1fbc700000000,
104'h08b5a5306b072b2d0e00000001,
104'hb819a8333347ca558f00000000,
104'hbc165c252cb860a87000000000,
104'h9435b05b6b4c88bd9900000000,
104'h94f54edaea4b14db9600000000,
104'h54070f350e9f6c6c3e00000000,
104'h54969c602debc05ad700000000,
104'h9ce645aacc97ae642f8604200c,
104'h34b3b2826776ab87edffffffff,
104'hbc41f16983774d5dee00000000,
104'h94d119c8a2884a7a1000000000,
104'h666478dbc871c9d3e300000000,
104'h282f01835e3959137200000000,
104'hb882772e04b4a2026900000000,
104'h28e08bbcc1a2b6e84500000000,
104'h547de851fbed8de8db00000000,
104'h3455d93fab05035d0a00000000,
104'h308a14e8148a7b3e1400000000,
104'h6664d59bc92ff9875f00000000,
104'h909c3e6838af49845e3377ec66,
104'h669cc31639858c460b00000000,
104'hbc550af7aa9d45f43a00000000,
104'h667086c3e1b4c2346900000000,
104'h28ceb1829d0867891000000000,
104'h9083b468070851af108be5c717,
104'h287be5b7f7964afe2c00000000,
104'h34265a974ce4fcd0c900000000,
104'h340384010782eed20500000000,
104'h04cb8e9697d3ad76a700000000,
104'h9cc4fd8a89272f414e042d0008,
104'hb806b8750d33513b6600000000,
104'h30718441e3dd0244ba00000000,
104'h005b9effb76e757ddcca147d93,
104'h90e5f6d0cb7d739bfa98854b31,
104'h60ed33beda50a355a100000000,
104'h30318ca5637460bfe800000000,
104'h54d71f02aed77ba2ae00000000,
104'h2c7541e9ea25f4eb4b00000000,
104'h9cbe0bd47c9b92fe379a02d434,
104'hbc08038b1021e51d4300000000,
104'h94e2b400c5ad0dc65a00000000,
104'h000b9b3517606c13c06c0748d7,
104'h08c3ac14877ffc17ff00000001,
104'h085e5b55bc8506440a00000000,
104'h5419ef5b334475cb8800000000,
104'h94958b142be2edf0c500000000,
104'h60bc2bde78c6767c8c00000000,
104'h346c9261d9bf57127e00000000,
104'h30b4ce6e69b1798c6200000000,
104'hbcd4e5e6a90d6b651a00000000,
104'hb896ce942dd3d612a700000000,
104'h6092b31025a006664000000000,
104'h00dd3a9ebabddaee7b9b158d35,
104'h9c124c0b248d31501a00000000,
104'hb8e18394c3d8aab8b100000000,
104'h54e253c2c43f5f237e00000000,
104'h9cb4894869d0d7cea190814821,
104'h08fea9e2fd706895e000000001,
104'h94e66640ccf0c04ce100000000,
104'h66d816d8b00a48251400000000,
104'h3408fbcd11c6aa0c8d00000000,
104'h08c4b7ce89a9960e5300000000,
104'hb8793df9f2329eaf6500000000,
104'h90452ab18a3dc44f7b78eefef1,
104'hbcbb3f8e76b8078c7000000000,
104'h9c4a7a2d94031aa106021a2104,
104'h6074fe1be9af09c05e00000000,
104'h3068c9add1d2727ea400000000,
104'hb8d3ede8a7b1a2286300000000,
104'h60a2c15e4582b3280500000000,
104'h60e94606d2608163c100000000,
104'hb839ba2b73d80d96b000000000,
104'h08490c3f925ba7c7b700000001,
104'h30aea9c25d3cf8897900000000,
104'h60f7e11eef0ac1731500000000,
104'h04dfce8cbf40ec778100000000,
104'hb8738bf1e79142402200000000,
104'h54ef1bb8de98df9e3100000000,
104'h666246c1c40a41d11400000000,
104'h005d6533ba1d81fd3b7ae730f5,
104'h2834ca5d69e8177cd000000000,
104'h90864ba20c03394b068572e90a,
104'h9cc71a4e8e13b65f2703124e06,
104'h0868e879d147dd098f00000000,
104'h66cc10e49827c9554f00000000,
104'h086939e1d212326f2400000000,
104'h348fab281fe38efcc7ffffffff,
104'h04764ec5ec7f287dfe00000000,
104'h005c14e7b8b175ae620d8a961a,
104'h60c132d08218d3eb3100000000,
104'h288d74ac1add7788ba00000000,
104'h00f09a70e1f32b36e6e3c5a7c7,
104'hbc2077c540d73664ae00000000,
104'h087d4ed3fa2a829d5500000000,
104'h2c479e3b8f9bd7e23700000000,
104'hbca359e2463fc8197f00000000,
104'h545346dda623a15d4700000000,
104'h0013f249278e7f661ca271af43,
104'h08f87b34f06f53edde00000001,
104'h60542777a8d87e00b000000000,
104'h2cc27b90849148702200000000,
104'h94744d93e8a367264600000000,
104'h303b0af976ce4b849c00000000,
104'h288c298c18e3e7d0c700000000,
104'h90157b3f2ab2398664a742b94e,
104'h9427dd0f4f32b2bd6500000000,
104'h006878e9d0b45a8c681cd37638,
104'h2891928623873c680e00000000,
104'h08c2974685c77e788e00000001,
104'h28a3e91e4734370d6800000000,
104'h2ca59c644bf1d8e4e300000000,
104'h089120c222a1cea44300000001,
104'h94b48d0c69c89d2c9100000000,
104'h04cb06209601a4f10300000000,
104'h90a078ca406b5a6bd6cb22a196,
104'h54f79ea2eff88d6af100000000,
104'hb8a005ea405b177db600000000,
104'h289e94743dfa094cf400000000,
104'h2cfdbd7afb492eff9200000000,
104'h2cfb6284f6d18396a300000000,
104'h9c09174512b9eb4c7309034412,
104'h2c20407d40954d002a00000000,
104'hbc7645d7ec16e2832d00000000,
104'hbc55cecbabff5808fe00000000,
104'h2cf8c27af18d127c1a00000000,
104'h66638299c7e7b4eacf00000000,
104'h9ca4993c49d2bcd6a580981401,
104'h282cd1d3595ccda3b900000000,
104'h606274ebc4b102ea6200000000,
104'hb8cf1f269e9561ec2a00000000,
104'h90826b0e04ed41d8da6f2ad6de,
104'h602c65ff58b843427000000000,
104'h943987f773ee2e78dc00000000,
104'hbc8ea6861d35d0e56b00000000,
104'h54961aac2c38b1697100000000,
104'h04d011aca02f33cb5e00000000,
104'h6636c0fd6da083044100000000,
104'h9c33f51b67275ab34e23501346,
104'h30d03374a0c887689100000000,
104'h04dc673eb8f9b618f300000000,
104'h904dd15f9b4eea719d033b2e06,
104'h0888b34211d2b438a500000001,
104'h2c18ecc731c0fbb88100000000,
104'h6008851311a5fd0e4b00000000,
104'h54d2d67aa532ca9b6500000000,
104'hb88fd55c1f5e6e57bc00000000,
104'h288daa041b1682372d00000000,
104'hbcd7958aafc3d78c8700000000,
104'h9c4fd9b39faf85645f0f81201f,
104'h08b71bca6ed275eaa400000001,
104'h9c6e7a8fdc3d4ac37a2c4a8358,
104'h90a24f044400306f00a27f6b44,
104'h340a506514b9f8ac7300000000,
104'h543892eb71ab93d65700000000,
104'h04bb99c077c8c13e9100000000,
104'h2cd073e2a0b08e9a6100000000,
104'h66389bf1712ffe555f00000000,
104'hbcac131c58deecf8bd00000000,
104'h0482ef0005fb0d8af600000000,
104'h3442528384ce94ec9d00000000,
104'h60e789bacf1fec3b3f00000000,
104'h30c8c0c2914d82319b00000000,
104'hbcdd8daabb4493858900000000,
104'h04ea4546d4638245c700000000,
104'h908fd31c1f001441008fc75d1f,
104'h34568c3dada7b0624f00000000,
104'hbc9d351e3ab3730c6600000000,
104'h2896328e2c63b185c700000000,
104'hb85b9d7bb7d64444ac00000000,
104'h304fb1e99fc0b0688100000000,
104'h90a9d0be53530805a6fad8bbf5,
104'h60e90cb6d2fa198af400000000,
104'h301bfa35374f46299e00000000,
104'h60323a2764521727a400000000,
104'h660ef7eb1d7b6a4df600000000,
104'h048452240843cd398700000000,
104'h00ee66a8dcc65fca8cb4c67368,
104'h60817958022f557d5e00000000,
104'h00b96dfe7210edc321ca5bc193,
104'h54618d33c37b7b6df600000000,
104'h54924c38243cd30d7900000000,
104'h60778fdfefe93848d200000000,
104'h08e4a260c9b3a2466700000000,
104'h285bd447b794ef082900000000,
104'h086e8043dd415dcd8200000000,
104'h66e6ea16cde1686cc200000000,
104'h3038306d70ded3babd00000000,
104'h54e949bcd2488eed9100000000,
104'h9c46c4298dc7b9ec8f4680288d,
104'h544bc06197cdeac69b00000000,
104'h00955f822af889fef18de9811b,
104'h66049bf5098eddf61d00000000,
104'h08a1454842f01d4ae000000001,
104'h080d97211baca0365900000000,
104'h3494a304295108f1a2ffffffff,
104'h084685518d8bfb061700000000,
104'hb8dc1d04b8beb9c87d00000000,
104'h34f0beb0e126c59f4dffffffff,
104'h94b31a52661250712400000000,
104'h942f4c2f5eeb20fed600000000,
104'h34f2d0bae5c33d4486ffffffff,
104'h90b7d3746f6473dfc8d3a0aba7,
104'h543010cb601f9c613f00000000,
104'h30a042f040aa26bc5400000000,
104'h60f3d1cce7b051a06000000000,
104'h04f53dccea501fd5a000000000,
104'h309a7dcc34e4e4a0c900000000,
104'h668547f40a54ff23a900000000,
104'hb825fd994be31cbac600000000,
104'h940cb217194a1a639400000000,
104'h9c0e84bb1d165d0f2c06040b0c,
104'h04ae459c5cb1390e6200000000,
104'h2cde1d7ebcdac074b500000000,
104'h0864b0b3c94c10679800000000,
104'h0822f4f3455ff58bbf00000001,
104'h2cd8b246b1d97f62b200000000,
104'h300466e3089fdaac3f00000000,
104'h54c80602907c8ac1f900000000,
104'h3486c9d60d04d9f709ffffffff,
104'h2ce91054d2c918fe9200000000,
104'hbc49fb1f931c05453800000000,
104'h60f74a66ee326e556400000000,
104'h904eaac79d6ef233dd2058f440,
104'h04546e25a85768bfae00000000,
104'hb80e67971c61561bc200000000,
104'h546a623dd4687bfdd000000000,
104'h9cf26b20e4ae621c5ca2620044,
104'h04b9e61873a36d884600000000,
104'hbcf525aaeae1df10c300000000,
104'h9041fde583a0d09c41e12d79c2,
104'h28fa8a44f5e90994d200000000,
104'h90ac1e8e58ef4238de435cb686,
104'h9c2b1ab956972e042e030a0006,
104'h906919c3d238651570517cd6a2,
104'h005db395bbba047c7417b8122f,
104'h2caac9e855eb9daed700000000,
104'h545c1823b819ccd93300000000,
104'h08e67e30cc2a8e435500000001,
104'h288e3e6e1c812ab20200000000,
104'h2c4c2685987352cde600000000,
104'h00585b47b0a8c16a51011cb201,
104'h005e3f93bc447d0988a2bc9d44,
104'h6637ae356fa290184500000000,
104'h60967ec42cb6d0706d00000000,
104'h9c6a0d87d4210d9d42200d8540,
104'hbcc33e4886c8be449100000000,
104'h66ac324658b6048e6c00000000,
104'h2889a90613d7a17caf00000000,
104'h085ac441b5e52f4cca00000000,
104'h2838a6b17182bad60500000000,
104'h6002260304a693f24d00000000,
104'h94d887acb1f3eccee700000000,
104'h002900d752b4a05c69dda133bb,
104'h5423712b464a37a19400000000,
104'h00e190c8c3c2062484a396ed47,
104'h90d28916a5a1f54843737c5ee6,
104'h906db0a7db7356abe61ee60c3d,
104'h346be219d7f6d582ed00000000,
104'h5401a5fb03b85f067000000000,
104'h087d27a1fadb99cab700000000,
104'h2871ad11e3e14418c200000000,
104'hbcef09dadec3915a8700000000,
104'h665644f7ac8b5e781600000000,
104'h28dd69b0ba59d533b300000000,
104'hbcf33b78e641d6858300000000,
104'h902044cf4022440b440200c404,
104'h54ed791eda6e0059dc00000000,
104'h087161a1e2603e61c000000000,
104'h949b8d3837f377d0e600000000,
104'h66dabb54b5ff2270fe00000000,
104'h907cf9d3f993fc8627ef0555de,
104'h90d9add6b3f88836f12125e042,
104'h66243fb548f70ddaee00000000,
104'h3462e1cfc5743d6de800000000,
104'h309faa703ff146e4e200000000,
104'h60b2f8ae659e01923c00000000,
104'h942cdc4d59677a85ce00000000,
104'h6697f89c2fed01e2da00000000,
104'h08c31a5886e98f52d300000001,
104'h669f78883e591557b200000000,
104'h34c0585e80e11bacc2ffffffff,
104'h30558c1dabb9b8ac7300000000,
104'h00c504ec8aefc1aedfb4c69b69,
104'h9c806fc6004aca6195004a4000,
104'h048a954c15d94b34b200000000,
104'h9004f4b1091306af2617f21e2f,
104'h0040d18b811585d92b565764ac,
104'h60dfacc6bfa843925000000000,
104'h90bde0747be5defacb583e8eb0,
104'h005ed6b7bd8d6cc81aec437fd7,
104'h288d13941a8abfb21500000000,
104'h348909ea12263fcd4cffffffff,
104'h2ca8733850f4a8e0e900000000,
104'h285ca28fb9fcc7d8f900000000,
104'h00690a6bd20d0f1d1a761988ec,
104'h0053ed91a7d499eaa928877c50,
104'h54f9f2f6f372f6c5e500000000,
104'h045a149bb4c7d0c08f00000000,
104'h345a216bb4474ff58e00000000,
104'hb81cca1b3969c8d3d300000000,
104'h9cb8f11071651289ca20100040,
104'h3066b53bcdab9c5e5700000000,
104'h9cb96ff472211a1b42210a1042,
104'hb8ee9de6ddfe5f60fc00000000,
104'h2ce86ae4d06dc20bdb00000000,
104'h08c758cc8eef1b92de00000001,
104'h2871396be2fe4170fc00000000,
104'h905c7357b8388c757164ff22c9,
104'hbcdd49d4bac5c72c8b00000000,
104'h08a79fb04f069b3f0d00000001,
104'h666a6d2bd4ee55d6dc00000000,
104'h040ae0c915e79af0cf00000000,
104'h3043e33f87235fcd4600000000,
104'h9cfb7648f6a744424ea3444046,
104'h34aa269654cc232a98ffffffff,
104'hb869889fd30f71b31e00000000,
104'h00d57882aa91c5ca23673e4ccd,
104'h669094f4214a9b7d9500000000,
104'h301f2d0f3e4d314d9a00000000,
104'h049c99363964139dc800000000,
104'h90bdb7047b38af0b7185180f0a,
104'h34500013a02201cf4400000000,
104'h001f73f13e01441f0220b81040,
104'hbc964cf22c351f8d6a00000000,
104'h08b0381e6013cd672700000001,
104'h00af88045f7a3417f429bc1c53,
104'hbc959a9c2b41db818300000000,
104'hb8606a31c0c950649200000000,
104'h54ae01345c9a4ec43400000000,
104'hb8534929a68ecb361d00000000,
104'h66de6c74bc11b3512300000000,
104'h3495c3522b29fd0553ffffffff,
104'h667b03a7f6565cffac00000000,
104'h9cdf2bdebecdbc0c9bcd280c9a,
104'hbc5660d7acec436ed800000000,
104'h300bb6b9175e984bbd00000000,
104'hbcc39cd2876c9dfbd900000000,
104'h30f86488f08ad7781500000000,
104'h66971b242e853fbc0a00000000,
104'h2cabaebe571831173000000000,
104'h9cf2161ae413b3932712121224,
104'h2c76f387ed234a5d4600000000,
104'h6064eabfc978181bf000000000,
104'h607ca1cbf9ccf24a9900000000,
104'h9cb424dc68fbbbacf7b0208c60,
104'h00c725368e911d98225842ceb0,
104'h344c4b0398e77866ce00000000,
104'h54dc9236b943a2c58700000000,
104'h9c306a7b60a5d0224b20402240,
104'h287b11f9f66eb60bdd00000000,
104'h08ef6350de0cc8811900000001,
104'hb8ea0e68d48f25661e00000000,
104'h9cebf452d7ab86da57ab845257,
104'h2c0c1e2f186a5495d400000000,
104'h6603870b07b7ac4a6f00000000,
104'h941db0bd3b79f90ff300000000,
104'h345fbbc7bff671aeec00000000,
104'h60cc7a38982996155300000000,
104'h94feb58efdbd83a27b00000000,
104'h54139f932761b89fc300000000,
104'h283e26357ce79e84cf00000000,
104'h5408a275119cf36a3900000000,
104'h66751a3fea58ea6bb100000000,
104'h66850d4c0a829af60500000000,
104'h9c6884fdd16f1737de680435d0,
104'h2c58df45b1c3417a8600000000,
104'h30268c7b4d793883f200000000,
104'h3071b849e3b2f2f26500000000,
104'h28949582291361ab2600000000,
104'h0822c50745dd311eba00000000,
104'h54bc0fa0780201c90400000000,
104'h04796ae9f28eaf781d00000000,
104'h2ca2012044e8ffbad100000000,
104'h284ab41b9510cf3b2100000000,
104'h9c3553116afa961cf530121060,
104'h90657b8bca12db652577a0eeef,
104'hb89fdd3a3f79ef4bf300000000,
104'h9c1558e32a7d04affa1500a32a,
104'h5406322d0cad81605b00000000,
104'h66e24c90c4a91d965200000000,
104'h94822b30049d2a3a3a00000000,
104'h94392bbf72bd16587a00000000,
104'h2ce43452c8b80b747000000000,
104'h9468cc59d1a338f04600000000,
104'h948758600e3e26697c00000000,
104'h2c1ff10d3fdc251ab800000000,
104'h30440ce58809b8371300000000,
104'h6057f545af268c514d00000000,
104'hb84dbe2d9b1455b72800000000,
104'h0858392db0b8add27100000000,
104'hbc871b420ed3c786a700000000,
104'h903e4db37c8792980fb9df2b73,
104'h009921f2324aa60395e3c7f5c7,
104'h9c36e0816dd80960b010000020,
104'h66d8eacab168b547d100000000,
104'h90536805a61562a72a460aa28c,
104'h34c835149017012f2effffffff,
104'h9ca88f6851a9eca653a88c2051,
104'h08bcb2dc790bb9571700000001,
104'h3421629942552f5daa00000000,
104'h04fa14f0f441cd198300000000,
104'h2c333a43663be8857700000000,
104'h284ad6db95b047946000000000,
104'h605e67d1bcadc79a5b00000000,
104'h60e3cae8c79d6ba23a00000000,
104'h5427a1714f5ce9d9b900000000,
104'h941e66253ca98fe05300000000,
104'h08f62e0aec83163c0600000000,
104'h9055cc5bab6dbaabdb3876f070,
104'h5402d1510530b9856100000000,
104'h34f29c16e549fe1d93ffffffff,
104'h904377a986c1a2288382d58105,
104'h94717aa7e2bf94127f00000000,
104'h04ffa242ff337c676600000000,
104'h08f06016e072ba29e500000001,
104'h00799309f3da0e3ab453a144a7,
104'h048ea3301db04db86000000000,
104'h9cd838a8b0ad335e5a88300810,
104'h94abc580571327e32600000000,
104'h083dda8d7b2c99535900000000,
104'h90d0ff52a1a5397e4a75c62ceb,
104'h2cb784e26f953b502a00000000,
104'h60d18bb4a398672a3000000000,
104'hb8713495e2e49e52c900000000,
104'h286db471db732543e600000000,
104'h665ac34fb5e5cd16cb00000000,
104'h08849e14094cd3e39900000001,
104'hb829937d534414198800000000,
104'h00a0d3ea4175dae7eb16aed22c,
104'h3462fc4dc55f7d95be00000000,
104'h546b9401d7a785ea4f00000000,
104'h90db75aab65f0d87be84782d08,
104'h9c52db1fa597a0482f12800825,
104'hbcd6843eadbcbdaa7900000000,
104'hbc6e30d5dc8bd1201700000000,
104'h08b365786647397b8e00000001,
104'h546e336fdc48b74b9100000000,
104'h00d27b84a4555a37aa27d5bc4e,
104'h2822e3f74578c565f100000000,
104'h081f794d3ea762d64e00000000,
104'h08e4b238c966ddcbcd00000001,
104'h906c4e7dd831fc1b635db266bb,
104'h9cec48c2d8a8ae9851a8088050,
104'h3088d38211cef07a9d00000000,
104'h906518dfca14cdab2971d574e3,
104'h60c33586868fa8341f00000000,
104'hb8c6a6988d20949d4100000000,
104'h043d227b7a2d65455a00000000,
104'hbcc094be8181bcc80300000000,
104'h3041b50783d33f64a600000000,
104'h28c570da8aafbb4e5f00000000,
104'h30882096103de0157b00000000,
104'h34003f3b00a0dd064100000000,
104'hbc0f1d571eecfe8cd900000000,
104'hb840c6e981df228ebe00000000,
104'h54fd1434fae29bccc500000000,
104'h9c2a9db155d0dc42a1009c0001,
104'h66b10ada622bfe8d5700000000,
104'h28b2f42065d1063ea200000000,
104'h00f04fb6e0306f4b6020bf0240,
104'h00b921827273645fe62c85e258,
104'h30dce5f2b981b4420300000000,
104'h6045efe38b105e3f2000000000,
104'h2c20b17b41aa4d705400000000,
104'h08bda80e7b749b39e900000001,
104'h047962fdf23570916a00000000,
104'h0410dd9121505e6da000000000,
104'h9c9123e222ecc51cd980010000,
104'h54b7fab46fc2a2b28500000000,
104'h66d00258a007e0550f00000000,
104'h08058c890b1bf6a93700000001,
104'hbc921d4c24c981309300000000,
104'h941b4ed936b518aa6a00000000,
104'hbcee9068ddc68c6e8d00000000,
104'h008df82c1b7552d5ea034b0205,
104'h94fb201af6d2c88ca500000000,
104'h6683c5d407649703c900000000,
104'h0438a58d714f59c39e00000000,
104'h30d9c7dcb3655ad1ca00000000,
104'h94943aaa2856fe0dad00000000,
104'h089bed0c37f23398e400000001,
104'h902926235204092b082d2f085a,
104'h54dbcef6b77b327bf600000000,
104'h30af875e5fcc20969800000000,
104'h90b23de064bf004e7e0d3dae1a,
104'h6643c28b87adb78a5b00000000,
104'h00f78cdaef3bb9b37733468e66,
104'h54f2ac94e5ab4b065600000000,
104'h94fe9daefd938b022700000000,
104'h943677296cd05dc2a000000000,
104'h605eacebbd810c5a0200000000,
104'h08505cafa0bc343c7800000000,
104'hb897ddd82fb75d966e00000000,
104'h902b0c57566e50b1dc455ce68a,
104'h541e86853dca02509400000000,
104'h0831d60b63d0af1aa100000000,
104'hbc193bbd32f87de8f000000000,
104'h54489679913bc1377700000000,
104'h2cdd9d0abb79af77f300000000,
104'h9cd0630aa0f02a7ee0d0220aa0,
104'hb8f7e0bcefa2edda4500000000,
104'h9064f5efc9423c338426c9dc4d,
104'h08491fdd9206e3ad0d00000000,
104'hb8beda0c7df3314ae600000000,
104'h6088623610682b4bd000000000,
104'h00e65716ccf42a84e8da819bb4,
104'hb8326a59641baad13700000000,
104'h28a31d72468eea5c1d00000000,
104'h00b4418c6836b01b6deaf1a7d5,
104'h9cd4b250a9b0510e6090100020,
104'h545c83dfb9a4ccc24900000000,
104'h601f9b9d3fd09896a100000000,
104'h005f6c1dbe0172290260de46c0,
104'h941b4bff36b550b06a00000000,
104'h30f99fd0f3d14d64a200000000,
104'h2ceccee6d9091ad91200000000,
104'h607dbb47fb776357ee00000000,
104'h90fa3480f48526480a7f12c8fe,
104'hbcd89d8cb101ec970300000000,
104'h3422bdb745286c015000000000,
104'hb8d8746eb0aaf1825500000000,
104'h04a7c8344fb8aab87100000000,
104'hb842887585a8a6365100000000,
104'h2cb27a66648922ee1200000000,
104'h9c83c8ee07a9868e5381808e03,
104'hbc222f7b444312df8600000000,
104'h9c8817e8101832253008122010,
104'h9c0fa35d1f2bf285570ba20517,
104'h6604562b080308590600000000,
104'hbc30deb561256f9b4a00000000,
104'h2c3f2f477e4384438700000000,
104'h3009e2f5136329a1c600000000,
104'h0824a583494158c38200000001,
104'h609616422c922dd02400000000,
104'h34305def606d4c71da00000000,
104'h08d66f8eacee3324dc00000001,
104'h347aac55f54fd5ab9f00000000,
104'h66706283e080965a0100000000,
104'h08f45f42e8c7768c8e00000000,
104'h54498b8d938515ee0a00000000,
104'h009d4c023ad2d8f2a57024f4df,
104'hbccc1bd698b04e1c6000000000,
104'hbc419aa18302aa770500000000,
104'h0440054d80d3f4e0a700000000,
104'h5409d1eb136f3879de00000000,
104'h0864e69dc91cd5f73900000000,
104'h2ce9a36ad3cdcc109b00000000,
104'h0838b73171e68edacd00000000,
104'h94b9776e7201c61f0300000000,
104'h009733342ee10ac6c2783dfaf0,
104'hbc86b9000d457b3b8a00000000,
104'h601e07973c03beb90700000000,
104'h9c66e1edcdc6cfc28d46c1c08d,
104'h6081be00038aa56e1500000000,
104'h2cd946c0b25393d3a700000000,
104'h943f68e17ef8fb60f100000000,
104'h5483a2c607719f47e300000000,
104'h08570f61aeddbaccbb00000000,
104'h60d5640aaafeadb8fd00000000,
104'h287ad96df5d5d7aeab00000000,
104'hb8ddb75abb33fa896700000000,
104'h00defbb2bd083bc110e73773cd,
104'h9c605441c0a99cce5320144040,
104'hbc96639c2c1782832f00000000,
104'h54f5090aeab5a36a6b00000000,
104'h662823575045752d8a00000000,
104'h30be06c07c42f0f58500000000,
104'h00c99dce934446bf880de48e1b,
104'h3000ed3501fbd7caf700000000,
104'h606972afd2f18ff0e300000000,
104'h66ae96ec5d647609c800000000,
104'hbc772a65eef70b40ee00000000,
104'h08a5a5384b40d1898100000001,
104'h9013a21b270d10eb1a1eb2f03d,
104'h543bcc257762b3ebc500000000,
104'h081637bd2c5ad2ebb500000001,
104'h0859de7bb3bb46887600000000,
104'h9412b5f9253058fd6000000000,
104'h903699c76d4c6e7d987af7baf5,
104'h9c4c003998163c9b2c04001908,
104'h007c3255f855e8a5abd21afba3,
104'h663f7eab7eef2504de00000000,
104'h30649f33c9da259eb400000000,
104'h30354a376aa703324e00000000,
104'h0418a62b3156e5c3ad00000000,
104'h6601188f02ac0de45800000000,
104'h005da7cbbb4d952f9bab3cfb56,
104'h00dfe818bf2d7d935a0d65ac19,
104'h345e2b5dbcf767bcee00000000,
104'h901e6c053cdc087ab8c2647f84,
104'hbc192aed3241350d8200000000,
104'h28f4383ee8a81e985000000000,
104'h08c41f4888eb1478d600000001,
104'h34bfad6e7fb9e5a673ffffffff,
104'h042bcbfb5767b91bcf00000000,
104'h908ea5041d9ef5243d10502020,
104'h08dfcb50bfd78dd0af00000000,
104'h609fdd2c3f69d24bd300000000,
104'h90b4da54693b9139778f4b6d1e,
104'h9c4924d1923f2c197e09241112,
104'h60e9e4d2d3bbf1aa7700000000,
104'h946e479ddc8cd7461900000000,
104'h9cfbd158f79e69443c9a414034,
104'hbc74b9fde9e68a52cd00000000,
104'h54f40d30e84859e19000000000,
104'h5460051fc04459798800000000,
104'h60bdd8667b68a91fd100000000,
104'h9082f2ee051ef2b53d9c005b38,
104'h94ce51c89c255c594a00000000,
104'h34f17a14e2a599c24bffffffff,
104'h942b42e156e8f4a8d100000000,
104'h089f6a023e09e41d1300000001,
104'h669cabfc392b8aed5700000000,
104'h94d7d6deaf9d35023a00000000,
104'h949510242a53abc1a700000000,
104'h2c794599f23bf96d7700000000,
104'h041c812b398af3821500000000,
104'h602297db4542a4198500000000,
104'h2cca6b9494226a494400000000,
104'h663cb813790869851000000000,
104'hbc9a22b234e29ff4c500000000,
104'h048d056a1a9bbbe83700000000,
104'h28262c914c638821c700000000,
104'h2cbc7fce783c87417900000000,
104'h54964df82c4816299000000000,
104'h94ffb3ecffd02d4ca000000000,
104'h9c4c567798f99926f348102690,
104'h08cb672e964b41879600000001,
104'h341bac57373ed7f97d00000000,
104'h284203c184cd05289a00000000,
104'h549798a62fcaed3a9500000000,
104'h08c5c4908be8a332d100000001,
104'h30c45330889fe3483f00000000,
104'hbcdba148b7582c5db000000000,
104'h0036ce836de1103ec217dec22f,
104'hbc4afa57951553252a00000000,
104'h546f43e7de7131f9e200000000,
104'h282604e54c93e7c62700000000,
104'h28fa7f68f4784a13f000000000,
104'hbc26f6df4d9a143e3400000000,
104'h34a5ebd64bad39e65affffffff,
104'h948df2f21bf25848e400000000,
104'h66d25ebaa4ff1e94fe00000000,
104'h9c6bb48bd7f3455ee663040ac6,
104'h30b1a46263fa6cf4f400000000,
104'h0804fbd30998fac03100000000,
104'h04facbd8f505cda50b00000000,
104'h60bab9b875ac61665800000000,
104'hb86132e9c252b901a500000000,
104'h94a2fbe64534280f6800000000,
104'h60da5220b41dd3253b00000000,
104'h04be98ca7d2b7f355600000000,
104'h307e48cbfc9b07ec3600000000,
104'h66779b8fef3a95157500000000,
104'h308f28f21ea966f45200000000,
104'h2cd4701ea8ecd1aad900000000,
104'h34f30366e62abf9755ffffffff,
104'h608bcf2817a0d2b24100000000,
104'h042cb3b1599afcf23500000000,
104'h94e56a16ca2e27a95c00000000,
104'h949f6c1e3e4341e18600000000,
104'h5413571726fccdc6f900000000,
104'h28a901ba5224c4ff4900000000,
104'h34703d11e00a6c0b1400000000,
104'h08def850bd776ca9ee00000001,
104'h30ce3fb69c194f333200000000,
104'h307a4e6df4582afbb000000000,
104'h00c2ab6e850525b70ac7d1258f,
104'h28be095c7c0319d10600000000,
104'h049a616834f97bd4f200000000,
104'h94e4812cc9b556c66a00000000,
104'h2863038fc605f7890b00000000,
104'h90df6ca6be129f3725cdf3919b,
104'h0034e08f694c548d9881351d01,
104'hb8f6ad56edaaac405500000000,
104'h2ca99fd253c420608800000000,
104'h9411db8923fa4ebcf400000000,
104'h2c2bad895750363fa000000000,
104'h5438924b71044b490800000000,
104'h948a669a14a1fb204300000000,
104'h34957b662a5df641bbffffffff,
104'hbcff04b4fe2659c54c00000000,
104'hb8081b6b104b8fc19700000000,
104'h348e4a421cf87ea6f0ffffffff,
104'h28115da122485fa59000000000,
104'hb872ee73e59654022c00000000,
104'h28a6e0164d1691892d00000000,
104'h54fcc930f9d2bdd4a500000000,
104'hbc38ff957132d0c76500000000,
104'h9c10bf25214195d98300950101,
104'h34f7a3aaef47a47f8fffffffff,
104'h00356dbf6a196789324ed5489c,
104'h2821caa543fc8b88f900000000,
104'h04d8972ab146ec258d00000000,
104'h9cebd58cd73cd8837928d08051,
104'h30394e53722e46a55c00000000,
104'h3448942f91d24dc8a400000000,
104'h0822e2e34555ffc9ab00000001,
104'h2ca1111842ef7976de00000000,
104'h54648d49c9f7c208ef00000000,
104'h34471d958e05d1690b00000000,
104'h9cb1daac6332d5a36530d0a061,
104'h662e9daf5d038f3b0700000000,
104'h0457d901af5c5c93b800000000,
104'h3039943573d54c46aa00000000,
104'h66f302ece6a94e925200000000,
104'h6022eeb145c75dac8e00000000,
104'h9011ebdd232e35235c3fdefe7f,
104'h90d41170a822f04545f6e135ed,
104'hbc70abfde1f0a77ae100000000,
104'h2cb1237e6222e4ad4500000000,
104'h34390c3b7286869a0d00000000,
104'h28281aa7501c6b413800000000,
104'h2c737241e67ef93bfd00000000,
104'h948e87761d77601dee00000000,
104'h94948c7c299127d82200000000,
104'h341a213934d2671ca400000000,
104'h34d3be18a74cb8b199ffffffff,
104'h008011f8006ec7ddddeed9d5dd,
104'hbcb64b006cc80bbe9000000000,
104'h948702840ec009b68000000000,
104'h9cfb43e2f68836be108802a210,
104'h0097e6662fbb4fca76533630a5,
104'h9cd43228a89ec12a3d94002828,
104'h301987eb334274f18400000000,
104'h9c1683ff2db920427210004220,
104'h2822d41f45c6e7c68d00000000,
104'h08d1b852a39df2fe3b00000000,
104'h60cfe6ce9f0046a90000000000,
104'h54764acfec53fe1da700000000,
104'h6645d6838b52bbb3a500000000,
104'h2c795fe1f2eee81add00000000,
104'h9431408b624118c18200000000,
104'h662130b342bdb5307b00000000,
104'h604b94f39706b36f0d00000000,
104'h54e63730cc57035bae00000000,
104'h28332283663501176a00000000,
104'h08951a082abf06587e00000001,
104'h54a1e2cc43f0f2d8e100000000,
104'h661d58a53aa343a44600000000,
104'h90cf06169e2c118d58e3179bc6,
104'h2cb8b73071680e79d000000000,
104'h34873f700ef559d0eaffffffff,
104'hb8d76a9aae83c3d40700000000,
104'h9047d0a58fbdd8007bfa08a5f4,
104'h54fd048efa63c671c700000000,
104'hb8685641d02d04395a00000000,
104'h347a1f75f4d73acaae00000000,
104'h2c1f538f3ee0de54c100000000,
104'h9caeca7c5dbb831e77aa821c55,
104'h30ed7e9ada35c9ef6b00000000,
104'h6041b59183667b69cc00000000,
104'h54bbcc3277f22a66e400000000,
104'h00781d5ff00a7565148292c504,
104'h66b83be07071bed5e300000000,
104'h049a7750340ff48d1f00000000,
104'h28bd63f27aacbe185900000000,
104'h0011dd9523212a21423307b665,
104'h00d0bd72a136b2cb6d07703e0e,
104'h04aa3b1254633119c600000000,
104'hbc03b02d071117492200000000,
104'h0025377d4a190a33323e41b07c,
104'hbcc35eae86edb1aedb00000000,
104'h0009e33913ac57ea58b63b236b,
104'h34633243c63cafd97900000000,
104'h005d2377bad7da7caf34fdf469,
104'h306e26f5dc2283614500000000,
104'h66aede225d6fabe5df00000000,
104'h080ad79315317da76200000001,
104'h9ca7e5e44f033bdf060321c406,
104'h2c7e49a7fc832bc20600000000,
104'h2804a62d09550be7aa00000000,
104'h0899797c328d72941a00000000,
104'h00a88f2651642b37c80cba5e19,
104'h089da6223bcf6ab49e00000001,
104'h083641bd6c8372ce0600000000,
104'h04e35d64c631fc816300000000,
104'h60587b9bb0ba81667500000000,
104'h045047cba0b83c147000000000,
104'h04a7c32c4f6c777dd800000000,
104'h9067b4a5cfdb854cb7bc31e978,
104'h54d8d3a0b100734d0000000000,
104'h3081e5fe03af57c25e00000000,
104'h049fc8e23f07ccd30f00000000,
104'h94761ca1eca8f2d65100000000,
104'h94740b9be81e11c93c00000000,
104'h9cc3641c86a6b1a04d82200004,
104'h0020fd3b417ec1affd9fbeeb3e,
104'h00041eb908932700269745b92e,
104'h90cf63e89e0cc9bf19c3aa5787,
104'h0038518570bff98e7ff84b13ef,
104'h30f39694e747c0f38f00000000,
104'h6032b04b65d47fa8a800000000,
104'h004c68e9986ae409d5b74cf36d,
104'h9c34699968ec1b6ad824090848,
104'h60ded752bdb1d17c6300000000,
104'h2883b2b8074056b18000000000,
104'h009a72fc347f058bfe19788832,
104'hb88913b6127abf15f500000000,
104'h30128dd325e0162ec000000000,
104'h30bf73607e8a81f61500000000,
104'h28782683f0abaf245700000000,
104'h0882e3400599c86e3300000001,
104'h90c0947681354de96af5d99feb,
104'h048a2ba4147ed35dfd00000000,
104'h94a4f3da4952bdb5a500000000,
104'h909717962ec4d7588953c0cea7,
104'hb8e6519ccc2f53875e00000000,
104'h2ca980e2532898c15100000000,
104'hbc0297670528ea1d5100000000,
104'h94c11c168224c7b14900000000,
104'h664637a78cb29dee6500000000,
104'hb8fa047cf4ea1c04d400000000,
104'h00e69986cdf9493af2dfe2c1bf,
104'h2c90082020df3156be00000000,
104'h289144f222c5bffc8b00000000,
104'h0814b3d1298423060800000000,
104'h2c9bce9837d8cbeeb100000000,
104'h30e41f16c855e82dab00000000,
104'hb8c083e281bce8907900000000,
104'hb8a47840480d6fa91a00000000,
104'h5413d6fd27c9bf1a9300000000,
104'h005c5057b8567c13acb2cc6b64,
104'h9c9e8ad43dd5628caa94028428,
104'h346ba72bd7da3fc8b400000000,
104'h9cc89f1491cf4b9e9ec80b1490,
104'h3073b743e739b8e77300000000,
104'h2880fc2a014114cf8200000000,
104'h66f981eef353cd47a700000000,
104'h34cddf409b70f659e1ffffffff,
104'h664f1b3b9ef32688e600000000,
104'h3432064364a202384400000000,
104'h040fb5f11fbfce067f00000000,
104'h00129bdf25ae202a5cc0bc0981,
104'hb83a6f9d741088db2100000000,
104'h3009e37f13f5c9a8eb00000000,
104'h2cb7dc8a6ff7f3e2ef00000000,
104'h08d2a550a56185f3c300000001,
104'hb8d653c8aca95fbc5200000000,
104'h04385a3d70f12600e200000000,
104'h9c08fb2111116cc12200680100,
104'h603817f57014c0932900000000,
104'h28f59320eb3e670d7c00000000,
104'h003e3cdf7ccb6e209609ab0012,
104'h089d03123af4627ae800000001,
104'h2c2cdc2b5943c4e98700000000,
104'h082aa503558916aa1200000000,
104'h0896e9c42d7a14e7f400000001,
104'h34b651be6ce37af6c6ffffffff,
104'h305c2655b81063d52000000000,
104'h2c052cd10a3b22797600000000,
104'h3091cb4a235c2933b800000000,
104'h041530872af3580ee600000000,
104'h3463f6d3c765ca39cb00000000,
104'h94ff79eafeadfa565b00000000,
104'h945bd7d7b755d5e7ab00000000,
104'h347d54c9fa7217a9e400000000,
104'h00369a036d8c00f418c29af785,
104'h541c07af38824a220400000000,
104'h943911c3725be1e1b700000000,
104'h04eb5fe6d63ed39f7d00000000,
104'h54ac2844582b6ce75600000000,
104'h6632fd7d652f79bd5e00000000,
104'h94ee0774dc6f3003de00000000,
104'h287a5f3ff41121d72200000000,
104'h344405fb88c04ef08000000000,
104'h2cefaeb6df832d060600000000,
104'hbc595349b2083f2b1000000000,
104'h28f94c32f2b0942a6100000000,
104'h041663852c7e43f1fc00000000,
104'h547e1abbfc10c3df2100000000,
104'h663d1b9f7af2aa3ae500000000,
104'h2c308c21611c38813800000000,
104'h66f5bd40eba3c4c64700000000,
104'h2ce86cead090da262100000000,
104'h903892d97198a81231a03acb40,
104'hbcd77068aea218b24400000000,
104'h28c05b90803da6577b00000000,
104'hbc247ca74830c7bf6100000000,
104'h90f17754e2be8b8e7d4ffcda9f,
104'h2c39b66f73e6baa6cd00000000,
104'h94e1d2d2c35a997bb500000000,
104'h08d14d4ca2d22084a400000001,
104'h046d9375dbae43945c00000000,
104'h008d078c1adca036b969a7c2d3,
104'h9004836709aeab165daa287154,
104'h66a48e3c493a34597400000000,
104'hb89c3d9638d2db00a500000000,
104'h2cf67926ecabc7465700000000,
104'h60f319aee6a6c40a4d00000000,
104'h28881ad810318f1d6300000000,
104'h080fd81d1fc3f8b28700000000,
104'h00400c9d808929b612c9365392,
104'h54aa0e0a54ec2934d800000000,
104'h54677a7fce9378b02600000000,
104'h9ce75164cec15f8c82c1510482,
104'h603e2f4d7c7e3d65fc00000000,
104'h609924d83257fb77af00000000,
104'h28ad60905a4d74f39a00000000,
104'h28e7a3d0cf9e6e6c3c00000000,
104'h66e53a98ca2074334000000000,
104'h3014ee792956b7afad00000000,
104'h28712c6fe24ec3c39d00000000,
104'h00c555be8a1da0353be2f5f3c5,
104'h280ef3df1d38bbff7100000000,
104'hbcf8474cf0bbb6bc7700000000,
104'hb8546977a867e103cf00000000,
104'h009df9903bbc0bc2785a0552b3,
104'h54f00c80e05afeabb500000000,
104'h0075d7b5eb04ad83097a8538f4,
104'h08104f09201a04933400000001,
104'h2ca1ada443ece3f8d900000000,
104'h603da1dd7b6da215db00000000,
104'h5419940f330d2ce11a00000000,
104'h30b340866656a251ad00000000,
104'h54ec9c5cd9c4f7b68900000000,
104'hbc02bd550521081f4200000000,
104'h94fa3cbcf43221b56400000000,
104'h2c8e4d501c2eea1d5d00000000,
104'h66907c16201631d92c00000000,
104'h3425d4474b570ea7ae00000000,
104'h2c1ade1d35e554e0ca00000000,
104'h54d2b0c2a57347d9e600000000,
104'hb8ce0f349cfb1944f600000000,
104'h349e48123c7a8f8ff5ffffffff,
104'hbcfc508ef8b0eb426100000000,
104'h2cdf5242be42e3658500000000,
104'h9c7ea415fdd250d6a4520014a4,
104'h9059e61db3c6e0b48d9f06a93e,
104'h905eb875bdaae5ba55f45dcfe8,
104'h043e452d7c8b209e1600000000,
104'hbcad95185baa176e5400000000,
104'h30d267bea47f53fbfe00000000,
104'h6033062f6658a12db100000000,
104'h045248e1a4771f67ee00000000,
104'h2c61c8a1c31bc7ef3700000000,
104'h9052f25da516b73f2d44456288,
104'h60bc761a780256730400000000,
104'h60b448c068cf3b9e9e00000000,
104'h009731082e9759342e2e8a3c5c,
104'h34ed9756db46d4638dffffffff,
104'h08e21098c4769a71ed00000001,
104'h9440dc2d81488d279100000000,
104'h28684cb7d01ede233d00000000,
104'h0420d40b4117f1452f00000000,
104'h00b02a0a603dde077bee0811db,
104'h28d5c680abc467dc8800000000,
104'h6667a605cf720597e400000000,
104'h302d11db5ad84fc6b000000000,
104'h9c09e2d1133dee137b09e21113,
104'h90bf77227e7fdba1ffc0ac8381,
104'h0029535952a99a7253d2edcba5,
104'h9c1a26253403adc70702240504,
104'h2c8aa74815cd73769a00000000,
104'h60d6896ead3334556600000000,
104'hbcfc770ef84303978600000000,
104'h666cd24bd91ac5273500000000,
104'h5497afd22f3773116e00000000,
104'h904d44c59a2179d9426c3d1cd8,
104'h28d4bf86a99bc3e03700000000,
104'h608c43aa186acbc5d500000000,
104'hb8a180d243aecdc05d00000000,
104'h9c2d1c875a17f00b2f0510030a,
104'hb863e723c7dcfa30b900000000,
104'h94d793a6afc4f3828900000000,
104'hbc956aa22ab1c0686300000000,
104'h66843014085d96cbbb00000000,
104'h28633441c656e169ad00000000,
104'h2c6b479dd625ea3f4b00000000,
104'h047f09a7fedd63e8ba00000000,
104'h9442cacd8592a9fa2500000000,
104'h080cf943194c50679800000001,
104'h5496d0ee2d4d59db9a00000000,
104'h2c59c63fb3312d1f6200000000,
104'h60c8e40e9180217a0000000000,
104'h66c614868c2e3a0d5c00000000,
104'h94020cfb044568358a00000000,
104'h2c1254c924c26cec8400000000,
104'h04239f3d47d73128ae00000000,
104'h60f7706eee472d398e00000000,
104'h9482c52005da372eb400000000,
104'h94b835a470dfd030bf00000000,
104'hbcfacbb4f5e0c8e4c100000000,
104'h341783592fd6d4ccad00000000,
104'h90a22ec4440164a702a34a6346,
104'h54df3534bea4dfca4900000000,
104'h282e64d95c1d14913a00000000,
104'h66e3cfa6c79d77a83a00000000,
104'hb8d26b40a4318a7f6300000000,
104'h2830ebd961fd809efb00000000,
104'h0024120948d2fc0ca5f70e15ed,
104'hb8ca63b694d778a8ae00000000,
104'h545407f9a8a9be945300000000,
104'h902e3def5c19738732374e686e,
104'h04c4a6a2898fa3361f00000000,
104'h608359ea06a8d6b25100000000,
104'h30cb7e4c96a912ca5200000000,
104'h0420dbd7414fd5679f00000000,
104'h9029a2075395e9ee2bbc4be978,
104'h66da58a0b4f8aca2f100000000,
104'h0886b39a0d9614fe2c00000001,
104'h663cc1f579729f1fe500000000,
104'h00faaf96f53dec177b389bae70,
104'h66a8123a50bcb1587900000000,
104'h60727945e4164f132c00000000,
104'h94f1b8a2e392258c2400000000,
104'h667b26b1f644818d8900000000,
104'h34fbc516f7b4b7b669ffffffff,
104'h34c00ca88015c6e52bffffffff,
104'h046cd445d93099936100000000,
104'h94478ab78f0abe331500000000,
104'h9c74bb97e9962e9a2c142a9228,
104'h9c3a972975be7e567c3a160074,
104'h3449f53b93e5880ecb00000000,
104'h2cc30b0886c571e88a00000000,
104'h30cbcc1897a7a0e64f00000000,
104'h664cae23995ff347bf00000000,
104'h667547e3ea7159e1e200000000,
104'h003503056a9ca88c39d1ab91a3,
104'h2c8cd8fe19cc35789800000000,
104'hb8b5d2f86b469f978d00000000,
104'h043cc49d7940d3eb8100000000,
104'h90967a0a2cbb29fe762d53f45a,
104'h540050a900ff2f32fe00000000,
104'h28eff308df8379240600000000,
104'h0091afca2360970dc1f246d7e4,
104'h280fa37d1f4dfa219b00000000,
104'h6044ad73893f6cf57e00000000,
104'h0444e7b389a371d24600000000,
104'h547a19cdf4e0a024c100000000,
104'h2c255eb94a73d8d3e700000000,
104'h6097f5c22feae99cd500000000,
104'h9c93f65a2756f77fad12f65a25,
104'h00b25f0064a7c8144f5a2714b3,
104'h0496b7202d1cc1f33900000000,
104'h34d13bf2a28a3c0a14ffffffff,
104'hb8c7505a8e09740b1200000000,
104'h2c7ea7c7fdb743ba6e00000000,
104'hb8ea6414d4d96d60b200000000,
104'h080a1e69140c17211800000001,
104'h60f99316f368cd55d100000000,
104'h60ac688058de23f6bc00000000,
104'h60ac48f2589acefe3500000000,
104'h9c784781f070c9bde1704181e0,
104'h604b47ef96dce53eb900000000,
104'h30c3e18e87dcd5acb900000000,
104'h085af51bb56196adc300000001,
104'h5476ed9bede5bec0cb00000000,
104'hbc686441d0ef19a6de00000000,
104'h90699f4fd3f8a1b6f1913ef922,
104'h900523ef0addb048bbd893a7b1,
104'h60c053188050fd0ba100000000,
104'h9cbdc96e7ba1c46e43a1c06e43,
104'h34effa22dfff2cf8feffffffff,
104'hb8973ccc2efdc3b2fb00000000,
104'h28d74658ae4ca77d9900000000,
104'h085ec4d7bdb7bb746f00000000,
104'h2c18966931b9f8527300000000,
104'h54d8d316b16eb4cddd00000000,
104'h28a0a1bc41927cf62400000000,
104'h909a8fda35ebd09ad7715f40e2,
104'hbc05e4810bd1e0a2a300000000,
104'h281a262d340b23771600000000,
104'h002ccba359d75854ae0423f807,
104'h0841cfd9831851bf3000000000,
104'h045ca0cdb9229ecb4500000000,
104'h2c91a16c233aeb8f7500000000,
104'h34b1366c6216b07d2dffffffff,
104'hb89c1632384e88c39d00000000,
104'h609553ac2a7e47a9fc00000000,
104'hbc695c37d242a4f58500000000,
104'h08b1e078634e184b9c00000001,
104'h300d60471ade3b84bc00000000,
104'h307dd17ffbe0cc1cc100000000,
104'h607c99edf983238a0600000000,
104'h605ad429b5a8be9e5100000000,
104'h546b9777d74d2be79a00000000,
104'h90eabaa2d513790926f9c3abf3,
104'h30c549ec8aa8f7305100000000,
104'h6609a7db131aee5b3500000000,
104'hbc041121083e97c77d00000000,
104'hbc98fb7a31c0774c8000000000,
104'h60798799f3cbebc49700000000,
104'h6006fdf10d6d8e5ddb00000000,
104'h2c510ea5a24ab9059500000000,
104'h2c3f4c677ef64bc6ec00000000,
104'h94d91a50b27e8927fd00000000,
104'h607004c9e0b9a1867300000000,
104'hb85f3d67bec645848c00000000,
104'h30cfb1c49f1b57593600000000,
104'h60aaf57255cd93389b00000000,
104'h664ff6c59f53c6b7a700000000,
104'h04e336c0c679ef21f300000000,
104'h28e8fbf6d15156e1a200000000,
104'h286ab85fd52f89db5f00000000,
104'h54e99a42d327b8cf4f00000000,
104'h60ff0016fe49e3bf9300000000,
104'h9c78475bf048e3419148434190,
104'h34262e774c6428ebc800000000,
104'h6030c1a56183ceae0700000000,
104'h94b78ac86fcd4d389a00000000,
104'h308a7c501484f1560900000000,
104'h940acf191543e8498700000000,
104'h6673cb4be7547b35a800000000,
104'h2c1a343534d5d174ab00000000,
104'h004dcf3b9b0e52031c5c213eb7,
104'h9ca33da6467f7bd7fe23398646,
104'h603521916acfcd409f00000000,
104'h601245bd24e7124cce00000000,
104'h54434079869732262e00000000,
104'h90c4c980894f53759e8b9af517,
104'h0434badd6990efb42100000000,
104'h66ee74bedc9e2da63c00000000,
104'h60a01c68400e9aa31d00000000,
104'h342cee0559131b012600000000,
104'h08a999885323a96f4700000001,
104'hbc96629c2c093d5d1200000000,
104'h94df7b6abea3f0544700000000,
104'h04ced2929de13a5ac200000000,
104'h34ab4bfa56ffdd50ffffffffff,
104'hb8701cb5e0eed754dd00000000,
104'h6683c1e0073a741f7400000000,
104'h66d0ca8ca10655650c00000000,
104'h90cb6c8e96f50a38ea3e66b67c,
104'h60f59c68eb058d690b00000000,
104'h3008202b104cc2df9900000000,
104'hb839d5517374cbfde900000000,
104'h00df21a4be05cb090be4ecadc9,
104'h66fa4716f41b6d7f3600000000,
104'h600212a7044055758000000000,
104'h044f1e419e243a054800000000,
104'h94f89d9ef1b356a06600000000,
104'h34a06e1e402d81715bffffffff,
104'h2872e1b7e52900c55200000000,
104'h60a17cbc4260f75dc100000000,
104'h66909eda21b8ffdc7100000000,
104'h60fecee4fd6f4f25de00000000,
104'h304921b992fc75a8f800000000,
104'h66caf422950b97e31700000000,
104'h9cdfefbabf37b5a36f17a5a22f,
104'h007612c3ec42587584b86b3970,
104'h0812330d2435c1056b00000001,
104'h04dc33d2b8c86b769000000000,
104'h9468e69dd15182cfa300000000,
104'h66b64f1c6c1d9b453b00000000,
104'h66dbc214b7e8cbb8d100000000,
104'h007a172ff41efdfb3d99152b31,
104'h34b0e5e261350e416affffffff,
104'h9c748553e9651175ca640151c8,
104'h344547318a45daa38b00000000,
104'hb8ab25945689974e1300000000,
104'h0829dbeb53991ada3200000000,
104'h30d022c2a03130e36200000000,
104'h2cc186be838d0ea41a00000000,
104'h00551267aa74bb51e9c9cdb993,
104'h304bc31797a8077a5000000000,
104'h306880cfd1066b710c00000000,
104'h3408111f1071e49de300000000,
104'h546a3d05d42ea9e15d00000000,
104'h66de21c4bc5b4f03b600000000,
104'h602264d5447caefdf900000000,
104'h60b6c2b26deeb56add00000000,
104'h00c730cc8ec6dee08d8e0fad1b,
104'hbc718a57e34708518e00000000,
104'h2c9d80363bd6e568ad00000000,
104'hb82343db468835f01000000000,
104'h94c0251e80dd9230bb00000000,
104'h2c091b2b12d56646aa00000000,
104'h2859f053b38a74921400000000,
104'h945c88f5b900f70f0100000000,
104'h005e7d5dbc6337afc6c1b50d82,
104'h60f3fea2e7f237c4e400000000,
104'h9c8dbe8a1bb6be5c6d84be0809,
104'h905c5263b87ce5a3f920b7c041,
104'h2c4e48e79c47ff3b8f00000000,
104'h2cd6eb1cad2667a74c00000000,
104'h90aa603c548ca0a41926c0984d,
104'hbc68ac83d114ca8f2900000000,
104'h607bc319f71b54b73600000000,
104'h00e5a2facb237cd346091fce11,
104'h289236c824a5f54c4b00000000,
104'h94a56fb44ad9cab0b300000000,
104'h3060d359c19b60023600000000,
104'h304c749b98bf1a247e00000000,
104'h547e0f93fc4d12339a00000000,
104'h04d5c05aab48e6e99100000000,
104'h34028d03053484fd6900000000,
104'h90c9ba5e935e7e7dbc97c4232f,
104'h2892a3f425b449386800000000,
104'h044d8ed59b2e7c1b5c00000000,
104'h089eaf763d70e385e100000001,
104'h60775aa7eed204bca400000000,
104'h942619534c1d683d3a00000000,
104'h0013178126f9c320f30cdaa219,
104'h600926171257d77daf00000000,
104'h34c447ce88a0a3c241ffffffff,
104'hbcb5810c6bf13920e200000000,
104'hb83062bf608050de0000000000,
104'h60b9884273bd78c47a00000000,
104'h949e003c3cc36e708600000000,
104'h008a588014c701c28e515a42a2,
104'h3034c4f1693196356300000000,
104'hbc88995611821b3a0400000000,
104'h04ca0e4a94d113a4a200000000,
104'h60100911205c0405b800000000,
104'h66e65e76ccba60007400000000,
104'h601dc8b93bc1cebe8300000000,
104'hb86f885fdf995e403200000000,
104'h04d9681ab27afdc5f500000000,
104'h66239baf471857253000000000,
104'h940cb1c519f3df32e700000000,
104'hb8d090d4a130b5256100000000,
104'h04563701acd3a8e4a700000000,
104'h2cf4b4f8e91d807f3b00000000,
104'h9ca29bda45fa5476f4a2105244,
104'h9c33d60d676b9b2fd723920d47,
104'h9c38a32171c23b428400230000,
104'h30cd2eb89a63bcefc700000000,
104'hb863fa5dc72172694200000000,
104'h30fe1268fcca2f3e9400000000,
104'h348ac5dc1506e6c10dffffffff,
104'h66fd5948fab049566000000000,
104'h2c39ecab730f38e91e00000000,
104'hb8fb8c46f7d3ac36a700000000,
104'h30742493e86d593dda00000000,
104'h9053d10da7c73e968e94ef9b29,
104'hbc4fbe239fa2e3d84500000000,
104'h04d99608b3e1e8f4c300000000,
104'h66af30a45e643c99c800000000,
104'h28eefe64ddaf118c5e00000000,
104'h90a0662440c46b1888640d3cc8,
104'h2cd00e0ca05cd85bb900000000,
104'h30aec7705d84b6b20900000000,
104'h303e95af7d64131bc800000000,
104'h60340813682402874800000000,
104'h347adeb5f5660947cc00000000,
104'h2873b257e709e96d1300000000,
104'h2c35174b6afbf01ef700000000,
104'h340d734b1ae99a02d300000000,
104'h90e37e5ec6f4269ae81758c42e,
104'h9c1226bb243872a5701022a120,
104'h28a94f9a523931797200000000,
104'h30c7a32e8f545d6fa800000000,
104'h54ba6f6c745e7737bc00000000,
104'h08e745f6ceb5ec3c6b00000000,
104'h60e7d6fecf8ebc0c1d00000000,
104'h00e33f1ec64a34ab942d73ca5a,
104'h9cc0c03c81585df7b040403480,
104'h947e9d6ffdd06c12a000000000,
104'h9c7491d5e99350b42610109420,
104'h30c41a7888d74394ae00000000,
104'h90618b31c35cd9c1b93d52f07a,
104'h2827a6834fb604086c00000000,
104'h04fc307cf8e50c54ca00000000,
104'h345eb49dbd9d6a0c3a00000000,
104'h607b76a7f68a05701400000000,
104'hb83b4691769c41fc3800000000,
104'h0875af5beb7ce7cdf900000001,
104'h6695b8ec2b33c3f56700000000,
104'hb85a3501b4ec97e6d900000000,
104'h9c114efb22d7afd0af110ed022,
104'hb873d6c9e77237fbe400000000,
104'h30477ec78e76292bec00000000,
104'h04e0049cc03b64057600000000,
104'h9ca5fd1e4be35362c6a1510242,
104'hbca6bb2a4d2e2dc15c00000000,
104'h540b898d17c4ad908900000000,
104'hb8df2fdcbe02d8a90500000000,
104'h00ef7a5ede582e95b047a8f48e,
104'h908d3ce01a0f55fd1e82691d04,
104'h94a0089e403321076600000000,
104'h60a38d1e474080b58100000000,
104'h08e35c18c6d4bf44a900000000,
104'hbc568849ad7d198ffa00000000,
104'h9407575b0ea88f6a5100000000,
104'h28abfec4576e8307dd00000000,
104'h002c23af58d47f54a800a30400,
104'h00f395c2e76b3d59d65ed31cbd,
104'hb8557d21aaeec09cdd00000000,
104'h9493f32e27ff2280fe00000000,
104'hb88ebe7e1d7764a3ee00000000,
104'h5458a9b1b14d623b9a00000000,
104'h042dad535bb1b87e6300000000,
104'h282ce4b959483e039000000000,
104'h900005e900396111723964f872,
104'hb8eed472dd7a8513f500000000,
104'h08efc74edf6f36f1de00000001,
104'h60c7d9c88fded06abd00000000,
104'h546a3f51d499e27c3300000000,
104'h043572676a007ec30000000000,
104'h3495d6762b5637d1acffffffff,
104'h66aee4b85d627099c400000000,
104'h00229c1145b352c866d5eed9ab,
104'h0493abec27e78428cf00000000,
104'h9441922b831672ff2c00000000,
104'h90cea3ee9db8d16e71767280ec,
104'h2c0eb98d1dc297d28500000000,
104'h3059f567b3e5a624cb00000000,
104'h3479ddc9f39fdc5c3f00000000,
104'h9c8fc1c61fb941ca728941c212,
104'h547a2125f49e937c3d00000000,
104'h28f38f34e782519a0400000000,
104'h2c1848b130d223caa400000000,
104'h60e074a0c0482c8f9000000000,
104'h089bc836371fa3a53f00000001,
104'h904805b590a9cf6453e1cad1c3,
104'hb8e68e44cd1c35273800000000,
104'h086dfedfdbe29898c500000000,
104'h34cb90249777222deeffffffff,
104'h664cb14999b0c4666100000000,
104'hb8ec15e2d80bb8511700000000,
104'hb80e2edf1c99a8ca3300000000,
104'h5467c64dcf76e4f3ed00000000,
104'h90c6364e8cc7b1808f0187ce03,
104'h546b72edd6cc912a9900000000,
104'h9458df03b17e1c05fc00000000,
104'h906aa411d5c8bdd891a219c944,
104'h663a052774de7390bc00000000,
104'h548fe4c21f985f943000000000,
104'h2c7175a9e27bcd23f700000000,
104'h30afcece5f15fabd2b00000000,
104'h2c0fda331ff7c378ef00000000,
104'h04cad6c29515ff6d2b00000000,
104'hb800653300a5330a4a00000000,
104'h60e9d7e8d31ee5813d00000000,
104'h66e33dd2c6ecb616d900000000,
104'h94e1604cc2a908925200000000,
104'h2c5cabffb9eee098dd00000000,
104'h9447bcbd8fc244028400000000,
104'h280504650aa03c4a4000000000,
104'h54a9c4c253b14ee86200000000,
104'h66e5546eca5b04adb600000000,
104'h04ca66ac94f4d824e900000000,
104'h042cce4959a2a2f64500000000,
104'h3078f383f1ba624e7400000000,
104'h308af4e01594ea282900000000,
104'h544a2b1794a8dfc45100000000,
104'h305a87e1b54512fb8a00000000,
104'hbc4007ef809b0ea23600000000,
104'h66892fb612fc77eaf800000000,
104'h2c2c4b5b58a594c24b00000000,
104'h08e7e98ccf1d11353a00000001,
104'h2c59c967b384dbc40900000000,
104'h2c50334fa021b0d54300000000,
104'hb8c874dc904ead039d00000000,
104'h34c9f7aa93f7fe86efffffffff,
104'h04082b4910038d970700000000,
104'h289e3a0a3cb033c46000000000,
104'h007e40f7fc5bda5fb7da1b57b3,
104'h0802829d053e97cf7d00000001,
104'h00a1ccf443eca3f8d98e70ed1c,
104'h66c90a4892cabb9c9500000000,
104'h087ab50df5804abc0000000000,
104'hb841a6c183c875ee9000000000,
104'h006f79cdde3edac97dae54975b,
104'h0837766b6ed69f3cad00000000,
104'h302dc27f5b0227f70400000000,
104'h00b74c766e1f8dc53fd6da3bad,
104'h5439a92f73f1a9e6e300000000,
104'h280adcd115b751826e00000000,
104'h906fc6abdf4217f3842dd1585b,
104'hb814a8212933b0316700000000,
104'h9c85fe7c0bb4c5346984c43409,
104'h90f8a7d6f179e14ff381469902,
104'hb8570af3ae32bc8b6500000000,
104'h04bdba1e7b7e0a15fc00000000,
104'h2c84c916099f9c923f00000000,
104'h5453cde3a7707983e000000000,
104'h66bd44b47ac033a48000000000,
104'h082acecf5594a4502900000000,
104'h04ae845a5dd0dbdea100000000,
104'h6646514f8cbde0fc7b00000000,
104'h30751553ea27971b4f00000000,
104'h0879fe91f32de3c35b00000000,
104'h301157a922fdeaf8fb00000000,
104'h903ac0817550fa9fa16a3a1ed4,
104'h302f8a2b5f3e7cd37c00000000,
104'hbc30adc76194094c2800000000,
104'h344e96639df26dc2e400000000,
104'h9c75b5d5eb504547a0500545a0,
104'h94119c9f23aa76a65400000000,
104'h302d0cd15a88b1cc1100000000,
104'h28483fe790ffc41aff00000000,
104'h08df57aabef55bd6ea00000001,
104'h54f9b20cf308927d1100000000,
104'h28c7980c8f9856223000000000,
104'h907e7f97fc5c89e3b922f67445,
104'h60fcd864f9d8752eb000000000,
104'h2c751bd5ea04da2f0900000000,
104'h082497dd49ddcb32bb00000000,
104'hbc1d2cd33a7416fbe800000000,
104'h0019f66133abe42a57c5da8b8a,
104'h3465975bcb61d3a3c300000000,
104'h28b5a09e6b35c1d76b00000000,
104'hb8b94af87225ff414b00000000,
104'h28a27c00446797b1cf00000000,
104'h2856cdf9adf000b2e000000000,
104'h54eb12b2d6e246f2c400000000,
104'h2cbe89687df59294eb00000000,
104'h94abbfa257e49a9cc900000000,
104'h9483d51207755f43ea00000000,
104'h00159a7b2b9e43663cb3dde167,
104'h308cc38419295cd95200000000,
104'h30ae23a85ce893ced100000000,
104'h948cae081984e9320900000000,
104'h3477b057ef20fc114100000000,
104'h004580ab8bdaa5ecb520269840,
104'h546e9671dda146284200000000,
104'h60dbc638b74614618c00000000,
104'h008718a40e1191d32398aa7731,
104'h0049743d92f4f1aee93e65ec7b,
104'h3418125d309010882000000000,
104'h2cbb7704762c52af5800000000,
104'h665e63c5bc6a818bd500000000,
104'h6665fd9bcb257fff4a00000000,
104'h28851dca0ae56dd0ca00000000,
104'h281b85cb379e91fa3d00000000,
104'h305e6e19bc4d24199a00000000,
104'h2cb2a82265baccbe7500000000,
104'h00b94b1c724c74df9805bffc0a,
104'h0406a3ed0d8ebc261d00000000,
104'h30ffe000ff452e5f8a00000000,
104'h341eab353d740fcfe800000000,
104'h548ab8b0152658954c00000000,
104'h60c7eec88f0137110200000000,
104'h2cd4addaa9fc313cf800000000,
104'h90ae6a325c40bd0d81eed73fdd,
104'h547b90e9f735e7d36b00000000,
104'h9cc06fc08084649a0880648000,
104'h30b99808735d1991ba00000000,
104'hb868f47dd1f00458e000000000,
104'h2cc38a2287bb0d747600000000,
104'h34ec9c32d99822a230ffffffff,
104'hbc37aae96f27b03d4f00000000,
104'hbcf5856eebd05194a000000000,
104'h048966c012fe5060fc00000000,
104'hb819d57f33054b0b0a00000000,
104'h5415bedb2bf41a1ee800000000,
104'h94e9046ed23ecca17d00000000,
104'h664c7521984c53739800000000,
104'h60cbe908972533b14a00000000,
104'h2c19f84133a658164c00000000,
104'h54c384d88726d95b4d00000000,
104'h907e0fa5fc61558bc21f5a2e3e,
104'h30d2902aa5192e773200000000,
104'h90fb477af651c709a3aa807355,
104'h089dc60c3b7197a3e300000001,
104'h904b1cad9644b18b890fad261f,
104'h9c8ef0481df2093ae482000804,
104'hbc82e8e6058c9fce1900000000,
104'hbc86b36c0d65635bca00000000,
104'h90958e942b945e502801d0c403,
104'h60e91ac2d2c78dde8f00000000,
104'h30dde4e4bb33774d6600000000,
104'h9c90e45821f55462ea90444020,
104'h2c1de3c33b406ebf8000000000,
104'h30f58cf6ebc002408000000000,
104'h661e8fd73d9cbe623900000000,
104'hbc901c2c2000be990100000000,
104'h54dca690b9b691b26d00000000,
104'h944ab0479507a8430f00000000,
104'h00ee0a1cdc3c41ef782a4c0c54,
104'h9c86ca4e0d82b1dc0582804c05,
104'h348bed64177d920ffbffffffff,
104'h08065a110cb83dc27000000000,
104'h2c6dc015dbb6aad26d00000000,
104'h04c38a1a87b17a106200000000,
104'h2860da9bc140d6b38100000000,
104'h00834bb606b07ca26033c85866,
104'h3048ea1f9164fdedc900000000,
104'h00aea2f05d0e1f151cbcc20579,
104'h04f51c92ea4be27d9700000000,
104'hb8beb2967d5b9ac1b700000000,
104'h90f60c9eec481c1d90be10837c,
104'h2c4788338f63e4c7c700000000,
104'h08606dafc075d44deb00000001,
104'h9c6da813db68c9ffd1688813d1,
104'hbc2877ef506c4245d800000000,
104'h34525941a4b7cb066f00000000,
104'hbc82144c047ce705f900000000,
104'h00c2b1888572b83be53569c46a,
104'h0071c873e3bc8944792e51b85c,
104'h083561796a280db75000000000,
104'h667a62cff4d1f182a300000000,
104'h28e3405ac6970f562e00000000,
104'h9013668b264665fb8c550370aa,
104'h6686983a0dbba4b67700000000,
104'h66543793a8d3e6a8a700000000,
104'h940d31e71afdf530fb00000000,
104'h9c00069500ed2948da00000000,
104'hb84920e99221c3e54300000000,
104'hb8de7cfabc7b5555f600000000,
104'h046c4f8dd8518baba300000000,
104'h000d28f11a8d800c1b9aa8fd35,
104'h08dacae0b5615b21c200000001,
104'h54b5a9646b75e869eb00000000,
104'h309fceb03f2570a34a00000000,
104'hbc549a01a990f3262100000000,
104'h949191842378964df100000000,
104'h9c7d3f33fab1e6c46331260062,
104'h30efd0acdf4e3dfb9c00000000,
104'h28c5f2248bf1677ae200000000,
104'h00091c3512ec5d48d8f5797dea,
104'h34494cc39259b345b300000000,
104'hb832e2e5652909915200000000,
104'h00e815bad0ac9de25994b39d29,
104'h60203e4f4047d3f38f00000000,
104'h5437ec776f3f4ccf7e00000000,
104'h2c637eb9c6d2e546a500000000,
104'h34cab52295a7b3424fffffffff,
104'hbca677324c8bda2a1700000000,
104'h603ac4ad75b7ce3e6f00000000,
104'h04e58986cb505efba000000000,
104'h2827ccc14f02a07b0500000000,
104'h94b97242728e8bd21d00000000,
104'h041087c721e6ee74cd00000000,
104'h547bd4b1f7a5008e4a00000000,
104'h66b524ee6adbba68b700000000,
104'h66d286dca54ac0c99500000000,
104'h9c6e7423dc7a8053f56a0003d4,
104'h94ed9d94dbdacfe0b500000000,
104'h04a5d2104b8331ee0600000000,
104'h04843862081f8cef3f00000000,
104'h2859d423b3d5f2b6ab00000000,
104'h045c0d95b8f9ced2f300000000,
104'h665bb487b71e93eb3d00000000,
104'h90e7b634cfffc024ff18761030,
104'h08b17e2462add0825b00000000,
104'hbc47ba0f8fef7b42de00000000,
104'h3048f8af91bc493c7800000000,
104'h54ba5bb0749166482200000000,
104'h66e7548ace1340952600000000,
104'h904624658c664f13cc206b7640,
104'h000196e903d716c6aed8adafb1,
104'h282b3037563d473b7a00000000,
104'h00e9c5b4d3ef85cedfd94b83b2,
104'h346739f5ce8d40201a00000000,
104'h667cd397f9499d699300000000,
104'hbc586729b02e66dd5c00000000,
104'h303d4bff7aef7f10de00000000,
104'h944ad41f95cf404e9e00000000,
104'h2886bf180db1da006300000000,
104'h047cdfe5f941850f8300000000,
104'h5445edcf8bdf2738be00000000,
104'hb8e63846cc7abd7bf500000000,
104'h3061b5cdc344a5718900000000,
104'h90cda5cc9be49daec929386252,
104'h34c0bd7e81751527eaffffffff,
104'h9cf997c6f3592187b2590186b2,
104'h3497e0122f11349722ffffffff,
104'h940770410ee6689ccc00000000,
104'hbc6d5975da8dfbbc1b00000000,
104'h543590036b3652516c00000000,
104'h60fcb24cf9b498526900000000,
104'hb8ac229e5835d9bb6b00000000,
104'h34e76c0cced829d8b0ffffffff,
104'h0810aa5b215831bbb000000001,
104'h08de6cdabc7d3d89fa00000001,
104'h34f04c46e091a0e823ffffffff,
104'h94b02ba660ef0a5cde00000000,
104'h004cdc2d99e61da2cc32f9d065,
104'h30679c1bcffe6d12fc00000000,
104'h3458a89bb127aa054f00000000,
104'h9467daa5cfe6a426cd00000000,
104'h282d06db5a406feb8000000000,
104'h9430986f6113cbd52700000000,
104'h30079ef90f249cef4900000000,
104'h9c3747656e471a198e0702010e,
104'h605a77c3b447fe718f00000000,
104'h540106350254daafa900000000,
104'h66bac2c275335d896600000000,
104'h54694c49d2782b13f000000000,
104'h047a6847f4959b162b00000000,
104'h66c155cc82f8767ef000000000,
104'h28785359f0ec8bb2d900000000,
104'h54344faf689cb1f03900000000,
104'h94737dc5e6a193ba4300000000,
104'h9c9c4398382858275008400010,
104'h28ecbc18d936034b6c00000000,
104'h30b3c3f867de2598bc00000000,
104'h9c63499fc6db323eb643001e86,
104'hb85057f9a0c494848900000000,
104'h08781463f0925c302400000000,
104'h6011a785232818e75000000000,
104'h0843c93387b03c806000000000,
104'h94b1674a62971c782e00000000,
104'h66eb9f98d7606a47c000000000,
104'h60e004b4c053babba700000000,
104'h0840e5e3818474620800000000,
104'h305a11efb4f73ce4ee00000000,
104'h08f74d18ee0abd6d1500000001,
104'h54a271e644c355f68600000000,
104'hb8bdf50c7b9917c23200000000,
104'h348d44461add1ea8baffffffff,
104'h9c4738458e2721814e0720010e,
104'hbc87917c0f6dd179db00000000,
104'h080b381116e46080c800000000,
104'h0447b6b38f6546a3ca00000000,
104'hb851287da2861e620c00000000,
104'h305291d5a55a3023b400000000,
104'h66cb5c5296d90480b200000000,
104'hbc816d9002c415b48800000000,
104'h28d2111ea43277f56400000000,
104'h5474ad51e98b10d21600000000,
104'h2c08fb2d111db59d3b00000000,
104'h949f39423ea948bc5200000000,
104'hbcfb918af760ae17c100000000,
104'h3456aa4fad5a2e6bb400000000,
104'h08fc1a02f834a1bb6900000001,
104'h041436272813789d2600000000,
104'h30517523a24e7ca79c00000000,
104'h9cd25b30a443dfcb87425b0084,
104'hb87faa35ff12f2b52500000000,
104'h66334c9d66939a322700000000,
104'h9c3733456e125b852412130524,
104'h90dc1e56b82297d145fe8987fd,
104'h043709216ea84e705000000000,
104'h2c30b10761007e5f0000000000,
104'h042d6f535a5afe93b500000000,
104'h9c5c5e1db8da655cb458441cb0,
104'h28638029c75656c9ac00000000,
104'h045363c5a69a52023400000000,
104'h04bf78ac7e1ed5b13d00000000,
104'h9c3910e972747351e830104160,
104'h6669c4abd35829a3b000000000,
104'h9456b135ad9e1dfe3c00000000,
104'h3020cab1413b8cbd7700000000,
104'h9c8f39141eaa888a558a080014,
104'hb80778090e19e0d93300000000,
104'h2cfbb1b6f74947319200000000,
104'h607a8cbff5058b970b00000000,
104'hb81c650738e287ecc500000000,
104'h9438a7a1718012500000000000,
104'h9ccac9ac954d0e7b9a48082890,
104'h90e91238d2c776208e2e64185c,
104'h34d82f1ab099f05433ffffffff,
104'h60cd4cd49a1f4fe53e00000000,
104'h080529770ab210ba6400000000,
104'h2c295a7d5231ac396300000000,
104'h04bdbdb07b415ca58200000000,
104'h54aecd025d63a77bc700000000,
104'h60c64d728c2bc6d15700000000,
104'h9cf690ecedb9c9c073b080c061,
104'h9cc5432a8a8803bc1080032800,
104'h30d5798aaaa822ec5000000000,
104'h54557e03aadc05a0b800000000,
104'hb8178ce92fea2698d400000000,
104'hb80d7de71a1738792e00000000,
104'h54ee0fd0dc3e48217c00000000,
104'h08a74f844e867e040c00000000,
104'h2c1c51cf38a1569e4200000000,
104'h543538476abde9be7b00000000,
104'h04af392e5e6598f1cb00000000,
104'h340f22591e343ce16800000000,
104'hb8cb8efe9741a9b38300000000,
104'h04e4c8a8c90c226b1800000000,
104'h2cdf0b08be3313416600000000,
104'h6620a2e141472b158e00000000,
104'h94401fdb80d0abb6a100000000,
104'h6087916e0f5e895dbd00000000,
104'h340886bf1168b0f1d100000000,
104'h60c1497c82fd8d7efb00000000,
104'h30b68bc06d06a48b0d00000000,
104'h283580f76b59e177b300000000,
104'h00e119aec23ce7df791e018e3b,
104'h0469da8bd3658501cb00000000,
104'h940a8613154e180d9c00000000,
104'h2ccc91a299d68996ad00000000,
104'h305e1d3bbc1229ed2400000000,
104'h9c97e66a2fc08e788180866801,
104'h2ce46e30c8b3461c6600000000,
104'h003a49d1743bfc9f77764670eb,
104'h347a56c1f41e64f93c00000000,
104'h086f497fde5702c7ae00000000,
104'h3496cf782dc3aa9c87ffffffff,
104'h28f53be2ea4c516d9800000000,
104'h30ab77a2560282e50500000000,
104'h2c8bac2617bb96cc7700000000,
104'h66abe14a575d7d6dba00000000,
104'h30a686364d5fbae3bf00000000,
104'h9c079d3f0f51e98fa301890f03,
104'hbc0202c1047edb6bfd00000000,
104'hbc230709466f326bde00000000,
104'h9403532f061007e12000000000,
104'h301ad0f73509fad91300000000,
104'h66920dae2452bd7fa500000000,
104'h545e5013bca6f9764d00000000,
104'h54d65928ac542343a800000000,
104'h006c8829d9f994a0f3661ccacc,
104'h0807d94f0f9e05ea3c00000000,
104'h66bff7c47f123e732400000000,
104'h9c395a87720b93ef1709128712,
104'h34b524346a1890c931ffffffff,
104'h60cd3e009a7fd98dff00000000,
104'h94f7e584efad293e5a00000000,
104'h60fea5a6fdf9fcc0f300000000,
104'hb8c3727e86cf452e9e00000000,
104'h00ab60265643394586ee996bdc,
104'h9c012caf02e21db8c4000ca800,
104'hbc4a94eb95329c996500000000,
104'h66122c61242e03b55c00000000,
104'h2cbc3020784281f78500000000,
104'h2ccf8ca29ff93bc0f200000000,
104'h345d0eb3baf3ce58e700000000,
104'h000d773f1a149a392922117843,
104'h008bea4c173aec7d75c6d6c98c,
104'hb8acf0c25977df39ef00000000,
104'h048b055a16f288dee500000000,
104'h000864791049d29d93523716a3,
104'h906a970bd5100dbb207a9ab0f5,
104'h9c46f06f8d702001e040200180,
104'h9c67f749cf15df0d2b05d7090b,
104'h66e2716cc482f2be0500000000,
104'h28ed8abcdbff5690fe00000000,
104'h006c4f03d8c051f6802ca0fa58,
104'h661f6ed73ea27fc04400000000,
104'h045d077dba5b3c81b600000000,
104'h2ca0e5c2414393dd8700000000,
104'h547a7be5f44284fb8500000000,
104'h9cfe826afdd635dcacd60048ac,
104'h0020fc07413b6dc1765c69c8b7,
104'h30e9147ad2286e815000000000,
104'h007b1271f6ec04eed8671760ce,
104'h902d54615af36840e6de3c21bc,
104'h9474106de83140616200000000,
104'h28144f45288deb5a1b00000000,
104'hbcf15a06e2dcd9b2b900000000,
104'h9098931831bc99ca79240ad248,
104'h289e720c3cb6ea3e6d00000000,
104'h289c1a8438dbeb4ab700000000,
104'h6657c609af5f4725be00000000,
104'h340af8f5155fe95bbf00000000,
104'h66003a49006a9d3dd500000000,
104'h5496c6942d65ab33cb00000000,
104'h344d75d79ad74d24ae00000000,
104'h0876cc53edd291d2a500000000,
104'h08d6ee7eadb607386c00000000,
104'h3458efd9b13d43f37a00000000,
104'hb873b4cfe7a227944400000000,
104'h086f5f95de9c6a103800000000,
104'hbcb300106665d215cb00000000,
104'h9046feb18d772a69ee31d4d863,
104'h90fb7a50f6e5ce54cb1eb4043d,
104'h54d29118a51364f72600000000,
104'h309d4c5c3a3123af6200000000,
104'h08d6a77aadddaf76bb00000001,
104'h90e2e9bec5507543a0b29cfd65,
104'h66a24b40440711630e00000000,
104'h2cec9cc2d9311de96200000000,
104'h34c06a9680147ffb28ffffffff,
104'h30e2d276c5c80c3e9000000000,
104'h2c0e046b1cdc1a36b800000000,
104'h9ccb26a696485ea1904806a090,
104'h08611467c22c24d55800000000,
104'h900c2fdb1809bf2b130590f00b,
104'h04ac3ef85817c6532f00000000,
104'h946c0b63d87a7fb9f400000000,
104'h944b3d4b96a582e84b00000000,
104'h0415a94b2b3975e77200000000,
104'h28e40948c85b7893b600000000,
104'h66f0d85ae133970f6700000000,
104'h9408c9a111e55b10ca00000000,
104'h04591225b2615451c200000000,
104'h28867dbc0cd02fdca000000000,
104'h04ff06eefe7fb685ff00000000,
104'h900c69c91817ca312f1ba3f837,
104'h5480e9c801e13a48c200000000,
104'h549842b23002070d0400000000,
104'h90057c7d0a326bf9643717846e,
104'h28d31a26a683c9280700000000,
104'h2ce5db98cbce43b09c00000000,
104'h604b0a8d962bb5035700000000,
104'h60320a6764fe414cfc00000000,
104'h2c35a3156b4eacd79d00000000,
104'h9c9c3ef2384248678400086200,
104'h902713a94ef20ca0e4d51f09aa,
104'h3416ee0b2d7c3c5ff800000000,
104'h2cea18f6d4afa61c5f00000000,
104'h60319739639b5c4c3600000000,
104'hb864a869c98f7cc41e00000000,
104'h040050cb00235f114600000000,
104'h34355c2d6a9341d82600000000,
104'h901a13cb34ab4f4256b15c8962,
104'hb8759f2beb6f9051df00000000,
104'h30f9c804f33027416000000000,
104'h08cc991499aee8ea5d00000000,
104'hbcce10069cd72d26ae00000000,
104'h66beda507d3a6e237400000000,
104'h0883d51a077c0ed1f800000001,
104'h04e6c80ecd0460350800000000,
104'hb897934c2f26bdd94d00000000,
104'h2c81c83a0350591da000000000,
104'h30f9656af2450b9f8a00000000,
104'h047e2d7dfcd54896aa00000000,
104'h540fd0ff1f44053b8800000000,
104'h54f5e344ebb5301e6a00000000,
104'h54a552544ae50f8cca00000000,
104'h28c1d9be83069eef0d00000000,
104'h904ca87b996ac32dd5266b564c,
104'h009231d4246bee07d7fe1fdbfb,
104'h2c87e13c0f798879f300000000,
104'h94b729326ef43c1ee800000000,
104'h04be25227c47f38d8f00000000,
104'h2c86c6440d4229b58400000000,
104'h90cc437c987ae045f5b6a3396d,
104'h940b443916b455046800000000,
104'h28bbfe5677c94e3a9200000000,
104'hb8663efbcc0b960b1700000000,
104'h94ee1678dc43fccf8700000000,
104'h94149f3329cafa809500000000,
104'h94c3177486dcc718b900000000,
104'h9cff4652fe4d81e79b4d00429a,
104'h668ee3901d89bff81300000000,
104'h28047a81084d99779b00000000,
104'h6662ffddc5200e074000000000,
104'hb86612adcc5a582bb400000000,
104'h94fba022f7c287a08500000000,
104'h0448628190767ac1ec00000000,
104'h66db72f0b6800ee20000000000,
104'h082de66b5bdd1fb4ba00000000,
104'h30622d91c47dada9fb00000000,
104'h041baf9537a843425000000000,
104'h0869d80fd3c8718c9000000000,
104'h2cd28feaa5d4fb66a900000000,
104'h00b6d9386dab07ee5661e126c3,
104'h0849061b92e173dcc200000000,
104'hb846c2998d2319e74600000000,
104'h2c51e98fa300aa210100000000,
104'h2849dc7d93d26854a400000000,
104'hb81bd673379fe96c3f00000000,
104'h345371efa687a7d00f00000000,
104'h30f559b4eaba06be7400000000,
104'h600cdcbb193b1cb97600000000,
104'h6081dcfe03345cd56800000000,
104'h3477516fee1af7293500000000,
104'h604b52bf964188278300000000,
104'h94886b5410036efd0600000000,
104'h605ca21fb985e2f20b00000000,
104'h34ad78785a7e9fcffdffffffff,
104'h0850d30ba179c135f300000001,
104'h348185a8032824ff50ffffffff,
104'h6602fa3105456ca78a00000000,
104'h28c22a6e841075a52000000000,
104'h9ccae4fa9512e0c92502e0c805,
104'hbc4f15199e7c00a1f800000000,
104'h54f28594e59146d22200000000,
104'h54c056ae801a088b3400000000,
104'h66d01eeca02631c54c00000000,
104'h00df6f02be8f3fc01e6eaec2dc,
104'h08b130ac62089a571100000001,
104'h940f189b1ef0245ee000000000,
104'h6082234204419b078300000000,
104'h666dd4c7db871c3e0e00000000,
104'h2cdeb3d8bd4eec119d00000000,
104'h943f37937e0251010400000000,
104'h04f7205aeee31f70c600000000,
104'hbce7f3c8cfe54bfeca00000000,
104'h94761377ecff9ce2ff00000000,
104'hb888a6f411da5252b400000000,
104'h54535097a6645de1c800000000,
104'h30036563063f80db7f00000000,
104'h903f1fe97e1169ab222e76425c,
104'h04f80620f00ba8351700000000,
104'h34127a5524561139ac00000000,
104'h2c032ef906e6e8b8cd00000000,
104'h906ff58ddfa9eb4a53c61ec78c,
104'hbc4c207998130e852600000000,
104'h04816ff6024b90599700000000,
104'hbc2d41eb5a7fad73ff00000000,
104'h9c7e7cc3fc6116a1c2601481c0,
104'h04836d5a0625fd234b00000000,
104'h04678fddcf164e1f2c00000000,
104'h66effb96df8874ee1000000000,
104'h9c21e9ed43f4bc8ce920a88c41,
104'h2c19902933f227f0e400000000,
104'h2ce04462c071596be200000000,
104'h04b7a55e6fd1e106a300000000,
104'h00843d6a086c09f1d8f0475be0,
104'h94f4d842e94cfecf9900000000,
104'h546483efc91cdd1f3900000000,
104'h0073f4a1e7e60fa0cc5a0442b3,
104'h9ca3c39a47ab07ac56a3038846,
104'h0003c10707d32d9aa6d6eea1ad,
104'h2c0450db0869a019d300000000,
104'h9ccd8abe9b601a97c0400a9680,
104'h60e494dcc9761a9fec00000000,
104'h008a71d414781c35f0028e0a04,
104'h54d0398ca034853b6900000000,
104'h9c0b7517163397cf6703150706,
104'h34d21592a4e583a8cbffffffff,
104'h08203e0f40056e7f0a00000000,
104'h5472d861e5520b63a400000000,
104'h90a8ad0a51e41922c84cb42899,
104'h6010761d2048dfa99100000000,
104'h665d2513ba8a84561500000000,
104'h90fa53b6f469cd73d3939ec527,
104'h2c9997f833acac785900000000,
104'h547e32d9fc7aa77ff500000000,
104'h903752436ebbf99e778cabdd19,
104'h94d1ddf0a342024b8400000000,
104'h2c41874183975baa2e00000000,
104'hb88594280ba3b00e4700000000,
104'h54109cff214326378600000000,
104'h34eb356cd67afcc7f5ffffffff,
104'h301838473084ac9e0900000000,
104'h089e2e6a3c6eaa33dd00000001,
104'h2c7408a5e8fd9dfcfb00000000,
104'h9c18248d30baabcc7518208c30,
104'h00ff5464fe23212f4622759444,
104'h90fe61fefcaba2ce5755c330ab,
104'h08834494062cb0d15900000001,
104'h289401ae28481a399000000000,
104'h2847f0ff8fd6b73ead00000000,
104'h547cdb47f96382c3c700000000,
104'hbc142c312894ea942900000000,
104'h54bd2f347a16eeeb2d00000000,
104'h2c680f75d09068ae2000000000,
104'h2ca212a2445b8eedb700000000,
104'h667e46d7fc8d93281b00000000,
104'h66fe9b7cfd42ecc58500000000,
104'h34601d25c095ab5c2b00000000,
104'h2ce9cc70d308e82f1100000000,
104'h301847e930002e6b0000000000,
104'h30e940e8d2fb72a4f600000000,
104'h04d07370a037f12b6f00000000,
104'h6634991169f40b66e800000000,
104'h9c658ec7cb57fc3baf458c038b,
104'h907da5d7fbdefb6cbda35ebb46,
104'h66bed7b67d7c27f7f800000000,
104'h606954e5d28c51741800000000,
104'h9cf3a6cee761787bc261204ac2,
104'h30a55ca84ac69dfa8d00000000,
104'hbc0bfb5917b239a26400000000,
104'h2c46a84d8d6b6f3bd600000000,
104'h08e7c760cf19db0b3300000001,
104'h60dc83bcb9018d310300000000,
104'hbc98fbb431fc8c0cf900000000,
104'h2c6487a7c908f5991100000000,
104'h003c53df786e97c9ddaaeba955,
104'hb80b4575160097ef0100000000,
104'h001ce22d39c781168fe46343c8,
104'h0865b355cbddd16cbb00000000,
104'h94ae5ba85cecde94d900000000,
104'h948f582e1e71a911e300000000,
104'h08aa241e5430f69f6100000001,
104'h545937b5b2f7cb98ef00000000,
104'h305b1a1bb6611b51c200000000,
104'h66757e4deacb477c9600000000,
104'h30e422eac85fc687bf00000000,
104'h9c4bed2797fd08fafa49082292,
104'h9c0d769b1a6675ddcc04749908,
104'h34e3062cc648160f90ffffffff,
104'h08e4abf4c9cb46ac9600000000,
104'h5409f80d139f8a723f00000000,
104'h903b848577e65216ccddd693bb,
104'h30af4a305e5253a7a400000000,
104'h60d17896a272c8f3e500000000,
104'h901048c72080ace40190e42321,
104'h04b403386887cfde0f00000000,
104'h002d30b95a5f5b27be8c8be118,
104'h5421ae3543051b370a00000000,
104'h60ae1bb25c84a92a0900000000,
104'h66fbde18f70f4b171e00000000,
104'h6024ac21493b236d7600000000,
104'hb8935e2e26f8075af000000000,
104'h90567931ac9614282cc06d1980,
104'h605bac85b7addb9e5b00000000,
104'h08fc3acef8c3bf5a8700000000,
104'h94d105e2a28fd33c1f00000000,
104'h9421b5a343d95ebeb200000000,
104'hbc9d31d83a40d5558100000000,
104'h6612671d2414ddcf2900000000,
104'h04c70eb28ed6c0bead00000000,
104'h667ef169fd5055cba000000000,
104'h9c78dd7bf18148180200481800,
104'h544747718e2349ab4600000000,
104'h08a94dfc52848dbe0900000000,
104'h941598e12beda22edb00000000,
104'h2cb34ac666237fcd4600000000,
104'h30b5fe266bc869ce9000000000,
104'hb8a8852251d5f41eab00000000,
104'hb8d6e46aad1848c93000000000,
104'hb8eac11cd5e68450cd00000000,
104'h289e399e3c3dc1197b00000000,
104'h6057e183af5429bda800000000,
104'h603f586b7e9f2a783e00000000,
104'h2c14b3df299399822700000000,
104'h9c7db43bfb086e691008242910,
104'h9cc27c7e848c607a1880607a00,
104'h04c8453a901c84213900000000,
104'hbcab426c56edbf42db00000000,
104'hbc59b459b354aca1a900000000,
104'h0030db7561b746366ee821abcf,
104'h0489473e12c96ea09200000000,
104'h348ab8241591317222ffffffff,
104'h28388c5b71c1529e8200000000,
104'hb89e6fc63c5084d3a100000000,
104'h5409c6d713c15ed68200000000,
104'h2c7f0c67fec2e7f28500000000,
104'h54cb1a9e969b53443600000000,
104'h54df16d2be9e422c3c00000000,
104'hbc42786184b5a5a46b00000000,
104'h60816294023016a16000000000,
104'h044649878c893d701200000000,
104'hb87499f9e928a0275100000000,
104'h66cedc3c9d10efe92100000000,
104'h04a58a0c4b9dad5c3b00000000,
104'h306c8f71d9a6bc044d00000000,
104'h66142e9d28213c9f4200000000,
104'hbc4ebecd9d8ac6821500000000,
104'h9cb77e306e87d8080f8758000e,
104'h60c76ebe8e1015e12000000000,
104'h28dbf618b7bab1767500000000,
104'h94f7b870ef2b0e575600000000,
104'hb888e66011b17e846200000000,
104'h0410f5cf21ddade0bb00000000,
104'h54387dd17070148de000000000,
104'h9056ad87adbd883e7beb25b9d6,
104'h30ee95fadda3c4ae4700000000,
104'h34cd3f029a8f82ea1fffffffff,
104'h007a3f25f43c77c378b6b6e96c,
104'h94414e6f82b5511e6a00000000,
104'h286e0c5fdc1d8a673b00000000,
104'h0413f0b927e8afdad100000000,
104'h341b1f7336c268f68400000000,
104'h04f7978cef8061d60000000000,
104'h949af4ee3572eb8fe500000000,
104'h0889bd52133aeb917500000001,
104'h28b3f01c6763720bc600000000,
104'h0475513bea4b0f459600000000,
104'h3424a70949dcc004b900000000,
104'h9c89e32e132208ef4400002e00,
104'hb8a1ee80434798dd8f00000000,
104'h08f38fdce7338a4b6700000001,
104'h9c93a60e27b81baa7090020a20,
104'h007facafffaf76d25e2f23825d,
104'hb85c4401b854df4fa900000000,
104'hb89a33d234ed5fc6da00000000,
104'h66b721606eb5ce606b00000000,
104'h946ff031df05c01f0b00000000,
104'h947985fbf316c33f2d00000000,
104'h3061697bc2d4f898a900000000,
104'h30c2745c84f9e404f300000000,
104'h34b2901665640bb1c8ffffffff,
104'h046535d1ca95be8e2b00000000,
104'h60232935467319a3e600000000,
104'h301aa663352b24775600000000,
104'h60dbfac0b7a19c6a4300000000,
104'h94c540e08a1ec71d3d00000000,
104'h00dcb762b97063c5e04d1b2899,
104'h2cd3ead4a7729399e500000000,
104'h00d6aa8aad19512d32effbb7df,
104'h668f808a1ffacecaf500000000,
104'hb820246540f8d3dcf100000000,
104'hb8df2110be6af14bd500000000,
104'h542ca5db590524d50a00000000,
104'h08cf3a329e1643772c00000001,
104'h9cb5cc986b8f42cc1e8540880a,
104'h28e75478ce00396b0000000000,
104'h9080ff0a0149ae4393c9514992,
104'h9c1a9f3335988f0231188f0231,
104'h286dd85fdb50e573a100000000,
104'h94df3c6cbe3f23d97e00000000,
104'h3039548172b1a0586300000000,
104'hbcb84cee706b974dd700000000,
104'h9421bc1943a8ccae5100000000,
104'h2c3ebc4b7d14a4772900000000,
104'h00575099ae9949f432f09a8de0,
104'hbc74ccc7e9b33e366600000000,
104'h34e5b826cb736565e6ffffffff,
104'hbcf06372e0fd6b24fa00000000,
104'h2c8229b2040a15f91400000000,
104'h282814195034e19f6900000000,
104'h666a58e7d491f86e2300000000,
104'h34eeed46dda563c04affffffff,
104'h0840223180460b438c00000001,
104'h34eb0446d6aedb665dffffffff,
104'h608df6ba1bee2ab0dc00000000,
104'h5492c1242577362bee00000000,
104'h28600871c0c34cb48600000000,
104'h66fceaaef920016d4000000000,
104'h081e36013ced7d0ada00000000,
104'h2c8f726e1e1bc6453700000000,
104'h9c92b6d42597992e2f92900425,
104'h005900b3b2ff2592fe582646b0,
104'h04c987189354cc5ba900000000,
104'h9ca1408442e9b3eed3a1008442,
104'h2c3493bb6953cb8da700000000,
104'hb8fbebb0f76295b7c500000000,
104'hb840a665819bd1823700000000,
104'h08ea96c4d544db078900000001,
104'h2c4711858e4f5ab59e00000000,
104'h28d93d0ab2179bbb2f00000000,
104'h08881c4410b0a1606100000001,
104'h28018c8f03edd36cdb00000000,
104'h549a2e903463d983c700000000,
104'h5480f21e01a9fd7c5300000000,
104'h3479bd17f32b2cd55600000000,
104'h94ad65445a4171038200000000,
104'h3025f5414b1876d73000000000,
104'h3074f44fe95b7cdfb600000000,
104'h0876293becf0c0c0e100000000,
104'h9c541045a86843a9d040000180,
104'h2c93fbf2273d7d937a00000000,
104'h902e98f95d0b57bf1625cf464b,
104'h9c464d138c4786058f4604018c,
104'h6617a8f12f76173dec00000000,
104'h08f8e508f1f7d494ef00000000,
104'h34d4217ca80dc7fd1bffffffff,
104'h902ce0ff595a017fb476e180ed,
104'h54a3f6a84779739ff200000000,
104'h60bddee07b3c7ebf7800000000,
104'h949e3b3e3cf3837ce700000000,
104'h6627e95d4f2a94115500000000,
104'h2cabecca577b1cb1f600000000,
104'h9cba23dc74bc1aee78b802cc70,
104'h00ed7f98da413c19822ebbb25c,
104'h0062368fc4f6fa98ed593128b1,
104'h04172ab72e6d9253db00000000,
104'hbc7c7a5bf83e64077c00000000,
104'h940ff3ef1f171fb72e00000000,
104'h34d4e4f2a90bcdf917ffffffff,
104'h30df7bcebe0c90631900000000,
104'h00c4b4bc896db0e7db3265a464,
104'h28b689a06dc858309000000000,
104'h2818dce93108030f1000000000,
104'h289e57703cac8ec05900000000,
104'h602d31635a12746d2400000000,
104'h341a9e0d35628b6dc500000000,
104'hbc6852d3d0906aba2000000000,
104'h00ca60fe94fa414ef4c4a24d88,
104'h54045aa908bebd787d00000000,
104'h94d37a94a6255b454a00000000,
104'h90d04710a07331dfe6a376cf46,
104'h94a4e7d849aa17ec5400000000,
104'h9c5626f5ace9b6ecd34026e480,
104'h005bd497b7e9e59ed345ba368a,
104'hbc920600243b615b7600000000,
104'h00d7675cae17be792fef25d5dd,
104'h942598a14b7b27a7f600000000,
104'h66474d758e7a4455f400000000,
104'h2cb4a80269345e0d6800000000,
104'h2cc106ea82d59cd2ab00000000,
104'h60d63e12acc6f2888d00000000,
104'hb827f28d4fd90d4cb200000000,
104'h28c691788ddd68d6ba00000000,
104'h047419e5e82c56dd5800000000,
104'h34c5b1a68bf89670f1ffffffff,
104'h0423bd414778d261f100000000,
104'h94cef2c29dcd1e969a00000000,
104'h00639fa9c78a4c7414edec1ddb,
104'h9c1519bd2aeeae40dd04080008,
104'h303a12ef7463a177c700000000,
104'h9c6f483fde04f82d0904482d08,
104'h54c0c39881e3197cc600000000,
104'h94a2a8b6458670d80c00000000,
104'h943944f772528469a500000000,
104'hb834da4f69b4ca7c6900000000,
104'h30885d1410ff15d4fe00000000,
104'h34331cf366573115ae00000000,
104'h946410bdc8b5011c6a00000000,
104'h001a3d51346e4661dc8883b310,
104'h28406f7b80bad55a7500000000,
104'h08cb40d296dddddabb00000001,
104'h34c71f9a8ea8996c51ffffffff,
104'h0838d1a571c878bc9000000000,
104'h0465aa2bcb36a7ef6d00000000,
104'hbc396ab5721882073100000000,
104'h943e86f57de04b3cc000000000,
104'h30aa43ac54734a71e600000000,
104'h3488e88611f61972ecffffffff,
104'h34cefcfa9d91c47823ffffffff,
104'h302b482b567c106df800000000,
104'h2c9a0bc834bb005a7600000000,
104'h301cb1ed39ef71c6de00000000,
104'h3049e60393dc6812b800000000,
104'h90d8d09ab1d05edaa0088e4011,
104'h9486ee560d7bbb5df700000000,
104'h08f2b9bee58b34c81600000000,
104'h2cee202edc7ecbb3fd00000000,
104'hb89279a6241da8693b00000000,
104'h66b47bb66884f8540900000000,
104'h30695f5dd293a2582700000000,
104'h28cf31dc9e4e6a3b9c00000000,
104'h9c6908add237daf56f2108a542,
104'h00cc904a996d1023da39a06e73,
104'h04492e25921436592800000000,
104'h3049ad6f933b5a897600000000,
104'h9ca82f0e501de0613b08200010,
104'hb8b0d47261d4b7a8a900000000,
104'h90525d77a42928a9527b75def6,
104'h54acb142598bcf7e1700000000,
104'h04fc0a2af8811e8a0200000000,
104'h947c3c8df81a7fc73400000000,
104'h287a50b5f4beed267d00000000,
104'hb81367bb268797fc0f00000000,
104'h6646a3638d3cf7557900000000,
104'h2cb488fa697e555bfc00000000,
104'h28d9173eb241b3b38300000000,
104'hbc6e8735dd939ede2700000000,
104'hbc2570154abe489c7c00000000,
104'h00abc61a57b501466a60c760c1,
104'h6646ec718d3ce82f7900000000,
104'h2cbdd2127bbd6b0a7a00000000,
104'h0026d1a14d5aec45b581bde702,
104'h0811cc4d23eba868d700000000,
104'h04a9b7b053eab27ad500000000,
104'h007996b3f3b69f5c6d30361060,
104'h2caf956a5f99382a3200000000,
104'h2cb5bff26b3b4ba17600000000,
104'h94f28c5ae5b376746600000000,
104'h902c2f7758407ab5806c55c2d8,
104'h2c9074cc20677e31ce00000000,
104'h2877916def8c47d21800000000,
104'h08cb29ce969d53fc3a00000000,
104'h9c3b82bf770757f50e0302b506,
104'h2c4b952b97438c358700000000,
104'h9c697d19d2e9d5d8d3695518d2,
104'h94f37b6ee6aba6f45700000000,
104'h54e282e6c5ee2dfadc00000000,
104'h900a07e514522c19a4582bfcb0,
104'hbc218b5743458a978b00000000,
104'h284f189b9e2e873d5d00000000,
104'h665aae55b5ca0fa89400000000,
104'h9c414a598266a3bbcd40021980,
104'h9c3b108976aad6ec552a108854,
104'h28a2c4ae450248b30400000000,
104'h94358f636b8dabdc1b00000000,
104'h6008c5e911fa34fcf400000000,
104'hb8082d0f10e287b8c500000000,
104'h0401ef1103befb367d00000000,
104'h08e63c76cce4cd78c900000000,
104'h541f4ff33e139dbd2700000000,
104'h30734d47e68645dc0c00000000,
104'h90ec331cd8d7eaaaaf3bd9b677,
104'h007ad7edf53fdb5d7fbab34b74,
104'h00a0a9d8411e97dd3dbf41b57e,
104'h2810a991218416360800000000,
104'h001ad83335ab1eee56c5f7218b,
104'h2c8610240c4f58679e00000000,
104'h346b00f9d6b3593a6600000000,
104'h665fc651bf11d9a72300000000,
104'h08fe51b4fc80dbe00100000000,
104'h66389f8171ef6376de00000000,
104'h04346eb5684e13b99c00000000,
104'h603cf3e17910cd0f2100000000,
104'h34ebbf02d77b2161f6ffffffff,
104'h9caacc5e5583376e0682044e04,
104'h9c50786ba0f67534ec507020a0,
104'h2882cea405e1094ec200000000,
104'h2cfa6b7af4752b51ea00000000,
104'h3055e921abc0ab2c8100000000,
104'h04258f7d4bd72790ae00000000,
104'h00dbbefcb7a503444a80c24101,
104'h54914e7c22d2f190a500000000,
104'h90bdd4247bebb192d75665b6ac,
104'hbc529149a5c550aa8a00000000,
104'h54c3794686f50bd2ea00000000,
104'hbca48b6a4940a7ff8100000000,
104'h284a77cd9481d97e0300000000,
104'h0084472e08b81264703c599278,
104'h28b87de27002cfd70500000000,
104'h08a2f1a245623e7bc400000001,
104'h9c514a77a255cdd3ab514853a2,
104'h28fae692f5300a9d6000000000,
104'h349d99323b2cd83159ffffffff,
104'h9c137c872672e0e7e512608724,
104'h904ece859d1ad56f35541beaa8,
104'h66bf90ce7f8ed3341d00000000,
104'h044b6397960209c50400000000,
104'h9ce2d376c5d47722a8c0532280,
104'h90501255a060532fc030417a60,
104'hbc89d346135e820bbd00000000,
104'hbc51c16da3b5256c6a00000000,
104'hb860c9d1c18f250c1e00000000,
104'h288c304818fd45f8fa00000000,
104'h0855275baa8929001200000000,
104'h28e96314d200480d0000000000,
104'h9ceddef4dbc0ca8481c0ca8481,
104'h542dcebf5bebc8a8d700000000,
104'h90a672684c8055f40026279c4c,
104'h341544f32a786a85f000000000,
104'h2858be45b1fc836cf900000000,
104'h664ca0199994921e2900000000,
104'h308185d2035492c9a900000000,
104'h04f42f60e850e1b3a100000000,
104'h66ebbf1ed79a27a23400000000,
104'h2816e2b52d8a753c1400000000,
104'h300e9ef71dbce55a7900000000,
104'h084236c3848ede781d00000000,
104'h2c2a64e554f5cb08eb00000000,
104'hbc2ae0f555b5e0e06b00000000,
104'h90efe736df0e4f8d1ce1a8bbc3,
104'h300a3b7914acedb45900000000,
104'h003edef77d9f3d7e3ede1c75bb,
104'h3420713740f05fece000000000,
104'hbc46f3f18d234f3d4600000000,
104'h948769e00eae78465c00000000,
104'hb81788b32f798ae3f300000000,
104'h004275dd8410193f20528f1ca4,
104'h006a4687d4335e4d669da4d53a,
104'h9036ba5b6da343104695f94b2b,
104'h5434697968ca7b149400000000,
104'h00785d47f0634fb9c6dbad01b6,
104'hb84acc57959a729a3400000000,
104'hb8187149309aeef23500000000,
104'h9424b4ab493a11f77400000000,
104'hb85fa1d1bf9be23a3700000000,
104'h90895ec012907e08201920c832,
104'h54219f0b430878cb1000000000,
104'h2cb449a668c20f688400000000,
104'h609549e02a2acba35500000000,
104'h943c432978d0ee74a100000000,
104'h54dd9ffebb95b97a2b00000000,
104'hb8c933ce928d6f481a00000000,
104'hb82f67d15e0ba2d11700000000,
104'h9c64aae9c9322dc1642028c140,
104'h903f9c857f66e5e1cd597964b2,
104'hbcf12a82e2c7e9768f00000000,
104'h00669a07cd001aa70066b4aecd,
104'h66143365282d21cb5a00000000,
104'h30a408fe48ce0edc9c00000000,
104'h2c9f11203e5d71d5ba00000000,
104'h346f8adfdf3b82037700000000,
104'h904265fd8454ac75a916c9882d,
104'h300225cd046ea153dd00000000,
104'h3418770930a9b8425300000000,
104'h288470b8087e43c7fc00000000,
104'h3052380fa4bd2b9c7a00000000,
104'h084d7f4d9ad0e61ca100000000,
104'h3413179d2617a89f2f00000000,
104'h901e8df73da166d042bfeb277f,
104'h08478afd8f53f925a700000001,
104'h04076de10e65821fcb00000000,
104'h34025a3b04b0eac86100000000,
104'h285fb0f7bf920e022400000000,
104'h08acac245926eaeb4d00000001,
104'h080095e701f8f638f100000000,
104'hb814d245299d62a23a00000000,
104'h30abb41a57bcf83c7900000000,
104'h3027d4e94f9bd2d03700000000,
104'h944a67bf94971f482e00000000,
104'h04e1bf1ac392b00c2500000000,
104'h3071fdc1e3ea005ad400000000,
104'h60c0aaa68197feb42f00000000,
104'h94589fcbb1deb630bd00000000,
104'h2cc68c1a8d33aee56700000000,
104'hbc27004b4e879d420f00000000,
104'h34d5bec0ab97b8782fffffffff,
104'h2c52c66ba5c4cfce8900000000,
104'h04f450a4e85ff70bbf00000000,
104'h286dba17db6661d1cc00000000,
104'h2cc20e9484b5c5fa6b00000000,
104'h0095affc2bc85d02905e0cfebb,
104'h942d501b5a735c61e600000000,
104'h30713587e2e47ce4c800000000,
104'h6032838565a2e91c4500000000,
104'h0864fce1c995aaae2b00000000,
104'h003279db64756ec7eaa7e8a34e,
104'h306e08f9dc8939601200000000,
104'hb82b72ef568d5fbc1a00000000,
104'h90cc99789919e1b333d578cbaa,
104'h66e0e946c138fa1b7100000000,
104'h346bd6cfd7107e232000000000,
104'h94be1e327cf863baf000000000,
104'h2cb23e24640686ed0d00000000,
104'h94ff65befe6b863dd700000000,
104'hbc26cd674de64e0ccc00000000,
104'h006e32b5dc83aafa07f1ddafe3,
104'h2c16ef432dc4fb3e8900000000,
104'h94bbe2a07794d70e2900000000,
104'h66292723521247fd2400000000,
104'h344749cf8ea2e7564500000000,
104'h94887d3410d9fb86b300000000,
104'hbcd8ff4cb1066c710c00000000,
104'h3014aa61299326d42600000000,
104'h04a268e4444546b58a00000000,
104'h30c3045886b920a67200000000,
104'h668b872417bb02407600000000,
104'h661c2983382a41755400000000,
104'h9c9b8156376cf2efd908804611,
104'h66826d0e04085f7d1000000000,
104'h9007f1870f26105f4c21e1d843,
104'hbcad02e85a970aba2e00000000,
104'h0436f0836db691ea6d00000000,
104'h6083ebb8075388e9a700000000,
104'h08bfe1d47ff34aace600000001,
104'h3448a0ef914291878500000000,
104'h9036ffcb6dd0c582a1e63a49cc,
104'h54b780b66f2fc9cd5f00000000,
104'h664fa76f9fb6210a6c00000000,
104'h048df9fa1b5b00bbb600000000,
104'h2ca1648c42e3ab9cc700000000,
104'h04a1786642cf2b089e00000000,
104'h281bbdb337893f561200000000,
104'h34731067e65f1f35be00000000,
104'h66f4c02ae9e85e12d000000000,
104'hb8ebeb28d704117b0800000000,
104'h349e4c003c9e0d703cffffffff,
104'h08ae72985c19cfd73300000001,
104'hbc0e20031cf072cae000000000,
104'h04283d5f50b4be046900000000,
104'hbc64a5bbc9bc2f3a7800000000,
104'h3050baeda10d917f1b00000000,
104'hbcbe7d767c5d7b9fba00000000,
104'h34c09f6881becd847dffffffff,
104'h08bcca3e79b104926200000000,
104'h2c8e0fc21c4fff0f9f00000000,
104'h30103de5200886751100000000,
104'h04198da5334ab8db9500000000,
104'h5412e4ef25af295a5e00000000,
104'hb8b7a37c6fd54f66aa00000000,
104'h043cb2ad79599d27b300000000,
104'h2ce35074c68f54ea1e00000000,
104'h60fecd2afd9df5723b00000000,
104'h30653479ca2bd5635700000000,
104'h34519933a34f459b9e00000000,
104'h089b7c363605528f0a00000001,
104'h300186510358fcb9b100000000,
104'hbcce8d189da77fe84e00000000,
104'h04869ad00d7601abec00000000,
104'h2c3e714b7c0abeab1500000000,
104'hb8f2bfc0e5df8f0cbf00000000,
104'h005503bbaafd59d4fa525d90a4,
104'hb842cceb85cfcf3a9f00000000,
104'h0828dc1351f6821eed00000000,
104'hb81e54dd3c743851e800000000,
104'h343cfac1794f0a079e00000000,
104'h60d230e0a4aba82a5700000000,
104'h542934ef529be1c83700000000,
104'h5411cd0323ac40645800000000,
104'h289760882ea653604c00000000,
104'hb8cb3410966d0259da00000000,
104'h90c1403c823dfe8b7bfcbeb7f9,
104'hb819db95336f2b27de00000000,
104'h605b2f75b6e094c0c100000000,
104'hb8242fdd48434fa78600000000,
104'h9c978e5c2ff35542e693044026,
104'h006fdff3dfe63876cc56186aab,
104'hbcaeede25d0a49091400000000,
104'h90f8e9a2f1d17df2a229945053,
104'hb818fbb131793ed1f200000000,
104'h2c17657b2e5be437b700000000,
104'h60622e35c42a87175500000000,
104'h9c0012c500c5771e8a00120400,
104'h344a309994777017ee00000000,
104'h306ba38dd70b66471600000000,
104'h54970ec82e7e81cdfd00000000,
104'h08b0c8a0615fa109bf00000001,
104'h00c92172923379f566fc9b67f8,
104'hb85cfd8bb9e03284c000000000,
104'h349bba003725080b4affffffff,
104'h2818149930ea5d92d400000000,
104'h90fe8ea0fdb44948684ac7e895,
104'h345e82d5bd2578d14a00000000,
104'h00f3e63ae73a04ad742deae85b,
104'h045e6c0bbc218a9b4300000000,
104'h007f8481ff55a6f5abd52b77aa,
104'h30036ec70625a50d4b00000000,
104'hb89255d82461fe99c300000000,
104'hb8fd3056fa8a02021400000000,
104'h549edb723dcbb7d69700000000,
104'h944ca8c799b9df187300000000,
104'h9442573984c598aa8b00000000,
104'h04a42ee048b919a87200000000,
104'h542eb7d95d967cce2c00000000,
104'h34a644304cc98ad293ffffffff,
104'hbc4144bd827d11c3fa00000000,
104'h2ccf21029e8c236e1800000000,
104'h9c720a13e4e552c0ca600200c0,
104'h669500642ab9c81a7300000000,
104'h080804c5106bc4c3d700000001,
104'h900b2c21164fed339f44c11289,
104'hbc3e0e7f7cea7286d400000000,
104'hb813c8c527ccf2d29900000000,
104'h344489ad898ba8881700000000,
104'h90ec619ad8d840d6b034214c68,
104'h284bcd7d979e71043c00000000,
104'h00a134b0427222dbe413578c26,
104'h080351db06a8cff65100000000,
104'hbcb33ece668764380e00000000,
104'h34b99b6e73f3bf1ae7ffffffff,
104'hbcfd0784fa84ac100900000000,
104'h6008e7a9118ce9ea1900000000,
104'h34a22d1e4445993b8bffffffff,
104'h00bc98b4797a29a7f436c25c6d,
104'h2c95b0a62b7b9e55f700000000,
104'hbc5b617db69ac1463500000000,
104'h080301e906689dbbd100000001,
104'h288231ac0472598be400000000,
104'h08a5cb724b8945881200000000,
104'h66fbe1b2f7d9bceab300000000,
104'h00dc7e8eb88b2b9a1667aa28ce,
104'h60419eb7835153a5a200000000,
104'h08019f4903aaa98c5500000000,
104'h90d016aaa0715fb5e2a1491f42,
104'hbc57d06faf5478b9a800000000,
104'h947d6437fab3f8d46700000000,
104'hbc949f8a29a70e3e4e00000000,
104'h00bbbac67794c8842950834aa0,
104'h66d610eaac2fb6f75f00000000,
104'h0874d287e9c285fc8500000000,
104'hb88eeb981dff737efe00000000,
104'h90ea1464d4de323cbc34265868,
104'h54b5c5606bf39432e700000000,
104'hb8c5860a8b0413fd0800000000,
104'h2c42ced185ce152e9c00000000,
104'hbc4775e78e1a73bb3400000000,
104'h54c85f329079ba4ff300000000,
104'h603ce72379a217b24400000000,
104'h04b240926495eb2e2b00000000,
104'h542abdab55847fe00800000000,
104'h9c77bbbfef264f294c260b294c,
104'h90d9aa2cb31be20137c2482d84,
104'h90cc64409802295d04ce4d1d9c,
104'h282ed6135d70e58de100000000,
104'h2c9ba464375f74a3be00000000,
104'h54fd4f88fa6a1fc5d400000000,
104'h345b0939b695bf982b00000000,
104'h303c357d78694fa1d200000000,
104'h30ff4e88fef4c89ae900000000,
104'h34cda3989b9259de24ffffffff,
104'hb8a02adc404ad9c59500000000,
104'hbcc25e4a84b804fc7000000000,
104'h6096db842d76e4f3ed00000000,
104'h54c63ebc8caa75325400000000,
104'h08a3708c46225fc14400000001,
104'h90215edb4263687dc64236a684,
104'h3464d8bdc97edf89fd00000000,
104'h907a0553f44c329b983637c86c,
104'h282fada75fa3756a4600000000,
104'h9043518f8699790632da2889b4,
104'h300fbf911fe5ca3ecb00000000,
104'h0084a7ba0978aefbf1fd56b5fa,
104'hb880618a004afaa39500000000,
104'h5465dcc5cb8b51761600000000,
104'hb827755f4eec32f2d800000000,
104'h94ac225858ebe332d700000000,
104'h609f379a3eeb0b4ad600000000,
104'h3413b2df27b8a8ac7100000000,
104'h001acb893551a387a36c6f10d8,
104'h2c323d8764e02420c000000000,
104'h34718735e3fa7f40f400000000,
104'hb84e123b9cab518a5600000000,
104'h30dcff6cb95c21d9b800000000,
104'h60560da9ac41a2a78300000000,
104'h2875d3bbebd46a66a800000000,
104'h28e6453acc22baef4500000000,
104'h043b3a6d76cfafca9f00000000,
104'h6605731f0a51eba3a300000000,
104'h9c314c8d62e79c9ccf210c8c42,
104'h9407223d0eaf6fba5e00000000,
104'h94e211e6c4d5cb3aab00000000,
104'h34be9a467dbb67f476ffffffff,
104'h2c4d4d099ad621c0ac00000000,
104'h60ee8ba2ddbe96cc7d00000000,
104'h5413073d26d4ee0aa900000000,
104'h54a17b804214dc7f2900000000,
104'h9464dc8fc984c1b20900000000,
104'h90d6efccad1573072ac39ccb87,
104'hbc0a07cd14380e197000000000,
104'h94b15b2e62d4ea20a900000000,
104'h60822e80041a80553500000000,
104'h2810c91721bce3487900000000,
104'hb812ecf725261d474c00000000,
104'hbc4649b18cb58db86b00000000,
104'h664c223d98f01d86e000000000,
104'h904c1de7985ce271b910ff9621,
104'hb84efc1f9d2989735300000000,
104'h90aea3645d87a0280f29034c52,
104'hbce3c324c76f9527df00000000,
104'h2c1200972408075f1000000000,
104'hbc2a669f54c7bc7e8f00000000,
104'h300090ab0176564fec00000000,
104'h0871c899e3e39f14c700000000,
104'hbc6e0f8ddc7704f5ee00000000,
104'h9081c9da03089c491189559312,
104'h601b85e537bac10a7500000000,
104'h946415f7c8372f336e00000000,
104'h34c7f5248fb42a1068ffffffff,
104'hbc77af33efee0ab2dc00000000,
104'h54d9c372b3bf4d407e00000000,
104'h905b3a9fb6a4f56049ffcfffff,
104'h28ece7bed936e1956d00000000,
104'h08fa0c04f4db659ab600000000,
104'h0071d5b3e3b343ca6625197e49,
104'h60c7f1f28f56dd7dad00000000,
104'h544929bd926f325fde00000000,
104'h94f7c1b2efed06e2da00000000,
104'h94081507108e498c1c00000000,
104'h9038a35171f58f66ebcd2c379a,
104'h2851897da3c13f508200000000,
104'h94461d9b8c3fc4697f00000000,
104'h907025cde083df6607f3faabe7,
104'h0456e21bad27ef014f00000000,
104'h001ce16139f0c74ae10da8ac1a,
104'h2836591f6c28700f5000000000,
104'h001e78653ce6e236cd055a9c09,
104'h3494edb029029c2b05ffffffff,
104'h902d97c75bfca528f9d132efa2,
104'h2cdb199cb65b57b3b600000000,
104'h9049c931937d0adffa34c3ee69,
104'h608b3170166772c3ce00000000,
104'hbc6b1f11d66a4fd1d400000000,
104'hb8fdf076fb03c5370700000000,
104'h2c3ca09179426e3d8400000000,
104'h6605c4bb0b550aa9aa00000000,
104'h004b759d96015a1f024ccfbc98,
104'h54c4db0a89cb7e789600000000,
104'h04d6d2e2ad9cfd303900000000,
104'h54c1eaf0832637bf4c00000000,
104'h082ca5cd59f6f2f2ed00000000,
104'h9407c2bb0fd2455aa400000000,
104'hbc3f00877e00049d0000000000,
104'h60db9370b7c189e48300000000,
104'h34de45febc89652e12ffffffff,
104'h6055fce5ab9557ba2a00000000,
104'h28c415de88ffad60ff00000000,
104'h94ead99cd5b8ccf87100000000,
104'h605af895b50b97b11700000000,
104'hbcabcae857c6ef788d00000000,
104'h28eecb4addd47c5aa800000000,
104'h08d184d4a35888dbb100000001,
104'h60b1ebec63608d5bc100000000,
104'h9cd7da2aaf15c2792b15c2282b,
104'h08c32528864ed26d9d00000001,
104'h3438887771a7816c4f00000000,
104'h66205a6940e6e50acd00000000,
104'h0490c40421e48294c900000000,
104'h3431f3db633a6c757400000000,
104'h28bd83e27b56368fac00000000,
104'h285b0a67b6d459a2a800000000,
104'h903a8ddb75f15db2e2cbd06997,
104'h2cba53be7431e3556300000000,
104'hbcd0427aa09e641e3c00000000,
104'h9c07ce490f0142030201420102,
104'h005c290db8ed7dacda49a6ba92,
104'hb83b2d3576e22beac400000000,
104'h04403b9d801281fd2500000000,
104'h9c67046fce2411094824000948,
104'hb8c4f2f8890488690900000000,
104'h66f4b49ee9be17167c00000000,
104'h2c7a12abf45d440bba00000000,
104'h2c2d17355a7cd595f900000000,
104'h30623501c4541fc1a800000000,
104'h60b9ea5c7321d1bb4300000000,
104'h94751705eaf11a28e200000000,
104'h948bfd0017f0ba88e100000000,
104'hbcc4a4828953619ba600000000,
104'h30521acda4e664b6cc00000000,
104'h0050c409a1a7b0344ff8743df0,
104'h666cb82dd99586c22b00000000,
104'h6655e2e1ab2a67d15400000000,
104'hbc0a5e4f146534e9ca00000000,
104'h90a2411644516e0fa2f32f19e6,
104'h04d8d71eb1ad1d245a00000000,
104'h903dfd797bf9c848f3c4353188,
104'hbc771945eeeb8332d700000000,
104'h2871e191e334f7996900000000,
104'h6693f4322710fc8d2100000000,
104'hb8f8edacf11214dd2400000000,
104'h28657c0fca9dec723b00000000,
104'h66e8a4d4d17eacb1fd00000000,
104'h94e535c8ca0dbfdd1b00000000,
104'h349c18da381b5b7336ffffffff,
104'h08fd030afacbe9889700000000,
104'h66adb6445ba029384000000000,
104'h0890ce4221ae9df45d00000001,
104'h54cbd062972ca5e55900000000,
104'h0410f69b21b34f586600000000,
104'h90f3ed40e79fc5103f6c2850d8,
104'h54017bff0278e9b1f100000000,
104'h6660d1a9c1d37a18a600000000,
104'h60a1eb1c43b3cebc6700000000,
104'h04374d276e581417b000000000,
104'h30a2095e449791f62f00000000,
104'h9cbdc6067b0b59e91609400012,
104'h088f40f01ef27498e400000001,
104'h90aa855655a7662a4e0de37c1b,
104'h9466ccc1cd76a1a3ed00000000,
104'h94d4c2e0a92543394a00000000,
104'h0078a479f16d29cddae5ce47cb,
104'h54547133a88f472e1e00000000,
104'hbc8728860ecebf949d00000000,
104'h30dcc996b99f2fe83e00000000,
104'h94cf8e149f7e3337fc00000000,
104'h30dd9818bb43ff038700000000,
104'h30670b0fce20aeaf4100000000,
104'h2cb747866eeb95d6d700000000,
104'h3018c22331cfb1b89f00000000,
104'h300dad6b1b2c11855800000000,
104'h90b06eba60a0cdce4110a37421,
104'h040596130b28e6e55100000000,
104'h945dd103bbbf22307e00000000,
104'h9cf91088f2cfbe949fc9108092,
104'hbc9cd9e8399297d62500000000,
104'h66ee7a98dcc910f09200000000,
104'h54ce97169d30dd7f6100000000,
104'h66de4cd0bcb882147100000000,
104'h666edefbdd1423a52800000000,
104'hb893a67a2728fddd5100000000,
104'hbc92bcbe25d39884a700000000,
104'h00b399a2674093e581f42d87e8,
104'h2c1b9c4f3759a41bb300000000,
104'h003737176e181387304f4a9e9e,
104'h08cb365896d3e422a700000001,
104'h66645a61c85267e3a400000000,
104'h28243c474858e819b100000000,
104'h341135cf224fb3d19f00000000,
104'h34c3c44687ffad36ffffffffff,
104'h28be9e6a7d182def3000000000,
104'h349f75403ee4da7ac9ffffffff,
104'h9cd51800aadabc98b5d01800a0,
104'h005472e7a859bca3b3ae2f8b5b,
104'h2810a11d219b51ea3600000000,
104'h3073099fe63902277200000000,
104'hb8e73f0cce6d07c1da00000000,
104'h2c731a99e61d37453a00000000,
104'h087649ddec53fbb7a700000000,
104'h66bd47be7af501f8ea00000000,
104'hb842785784aaeb265500000000,
104'h2cf4dfbee9311dfd6200000000,
104'h90d6ac06ada88f30517e2336fc,
104'h346e8a03dd8818d01000000000,
104'h540d7d391a60b8adc100000000,
104'h667fb2b9ff0bcdaf1700000000,
104'hb89186fa235d2c39ba00000000,
104'h0012b6cb250ca191191f585c3e,
104'h90e07316c0aa3e30544a4d2694,
104'h34abcfe457067f350cffffffff,
104'h66dcc61ab9f32eb0e600000000,
104'h04cac072959393162700000000,
104'hbcba6b50740a45951400000000,
104'hb8553fa3aa20c7734100000000,
104'hbcd200c6a4f8ae78f100000000,
104'h00762561ece00044c05625a6ac,
104'hbca6e3444d7214b7e400000000,
104'h301d56553a3417496800000000,
104'hbc2bfa5b5747ff6f8f00000000,
104'h600c6fef189297f82500000000,
104'h2c1344552638ed797100000000,
104'h081c345b38973b942e00000000,
104'h9cb4223c683731736e34203068,
104'h9026b6834dc525148ae39397c7,
104'hbcd463dea8038db90700000000,
104'h90c246128431dd3963f39b2be7,
104'h9c6013c9c0b790666f20104040,
104'h60b91b7872160e792c00000000,
104'h2cdc0344b89baf583700000000,
104'h54e9c3dcd30001130000000000,
104'hbc1f165f3e65242bca00000000,
104'h60fc4d30f823d7034700000000,
104'h9c9e4fe43cb788366f9608242c,
104'h2818321d300588030b00000000,
104'h9c579d61af86309c0c0610000c,
104'h6087060c0e789d93f100000000,
104'h082763214eb14a346200000000,
104'h08efe12cdfb1aeea6300000000,
104'h0814c82f29fab59cf500000000,
104'h94978c6a2fe59d0acb00000000,
104'h60e0c256c12ea3315d00000000,
104'h54d16d70a2b28eaa6500000000,
104'h9ce3e226c71bef0d3703e20407,
104'h348d32ac1a4eac499dffffffff,
104'hbc06dee90db83d0c7000000000,
104'h30ad3f485a389c217100000000,
104'h0461e2a9c38bd4cc1700000000,
104'h9091d73023e5be2ecb74691ee8,
104'h60ce96349d413da78200000000,
104'h90050b130aaa282e54af233d5e,
104'h3078ed17f1f49abae900000000,
104'hb8736459e6d6619aac00000000,
104'h283ab19b759ec6e03d00000000,
104'h001d512f3ac6dfb28de430e1c7,
104'h344dd0cf9bb830b67000000000,
104'hbcad50825a61416fc200000000,
104'h00a1667e42ef7698de90dd1720,
104'h9c5eddffbd3b4b8d761a498d34,
104'h94dd8932bb8fc2a21f00000000,
104'h66a21e104467a48bcf00000000,
104'h2ce1d63ac3f2e6b0e500000000,
104'hb8e849e2d0a450a04800000000,
104'h304abda3951b385f3600000000,
104'h6004db610966edcbcd00000000,
104'h60498e3393512d07a200000000,
104'h9c4f79399e02afc90502290904,
104'h34db417cb660b5c9c1ffffffff,
104'h3072a2d5e5e41c14c800000000,
104'h342a07c754d25b7ca400000000,
104'h34931c60269e85e83dffffffff,
104'h66a594204b3c1ac17800000000,
104'h2c3c1acb78474a458e00000000,
104'h041e28553c85fff00b00000000,
104'h543c2fbf785acbe1b500000000,
104'h9cee60f0dcbe83287dae00205c,
104'h085ef5a5bd272f3b4e00000000,
104'h94ffc13effdaa444b500000000,
104'hb8af7bac5e78d68ff100000000,
104'h6635ff4b6b7dc6dffb00000000,
104'h08af71c05e049dd90900000001,
104'h308d0fe21aa54e564a00000000,
104'h66af148e5ecbd6d49700000000,
104'h60f5f290ebd3f9c4a700000000,
104'h9c31d981637604fdec30008160,
104'hbcbe3da27c1900093200000000,
104'h040bdac5175c5991b800000000,
104'h2c0e6a231c0eebbb1d00000000,
104'h94a4034248c2ef888500000000,
104'h9ccadfdc95ae37385c8a171814
};

endmodule
