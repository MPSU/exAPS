`timescale 1ns / 1ps

module tb_rf_riscv();

    wire        CLK;
    wire [4:0]  A1;
    wire [4:0]  A2;
    wire [4:0]  A3;
    wire [31:0] WD3;
    wire        WE3;
    
    wire [31:0] RD1;
    wire [31:0] RD2;
    wire [31:0] RD1ref;
    wire [31:0] RD2ref;
    
    rf_riscv DUT(
        .clk(CLK),
        .A1 (A1 ),
        .A2 (A2 ),
        .A3 (A3 ),
        .WD3(WD3),
        .WE (WE3),
        .RD1(RD1),
        .RD2(RD2)
    );
    
    register_file_ref DUTref(
        .clk(CLK   ),
        .A1 (A1    ),
        .A2 (A2    ),
        .A3 (A3    ),
        .WD (WD3   ),
        .WE (WE3   ),
        .RD1(RD1ref),
        .RD2(RD2ref)
    );
    
    reg        clk;
    reg [4:0] a1;
    reg [4:0] a2;
    reg [4:0] a3;
    reg [31:0] WDr;
    reg        WEr;
    
    integer i, err_count = 0;
    
    assign CLK = clk;
    assign A1  = a1;
    assign A2  = a2;
    assign A3  = a3;
    assign WD3 = WDr;
    assign WE3 = WEr;
    
    parameter CLK_FREQ_MHz   = 100;
    parameter CLK_SEMI_PERIOD= 1e3/CLK_FREQ_MHz/2;
    
    parameter address_length = 32;

    initial clk <= 0;
    always #CLK_SEMI_PERIOD clk = ~clk;
    
    initial begin
      $display( "\nStart test: \n\n========================\nНАЖМИ НА КНОПКУ 'Run All'\n========================\n"); $stop();
      //------initial
      clk  <= 'b0;
      a1   <= 'b0;
      a2   <= 'b0;
      a3   <= 'b0;
      WDr  <= 'b0;
      WEr  <= 'b0;
      @(posedge clk);
      //----- reset
      for( i = 1; i < address_length; i = i + 1) begin
        @(posedge clk);
        a3  <= i;
        WDr <= 'b0;
        WEr <= 'b1;
      end
      @(posedge clk);
      a3  <= 'b0;
      WDr <= 'b1;
      WEr <= 'b1;
      @(posedge clk);
      WEr <= 'b0;
      a1  <= 'b0;
      @(posedge clk);
      if( RD1 !== 'b0 ) $stop("\n\nError of data with address 0\n\n");
      @(posedge clk);
      for( i = 1; i < address_length; i = i + 1) begin
        @(posedge clk);
        a3  <= i;
        WDr <= $urandom();
        WEr <= 'b1;
      end
      @(posedge clk);
      WEr <= 'b0;
      for( i = 0; i < address_length; i = i + 1) begin
        @(posedge clk);
        a1  <= i;
        a2  <= address_length - (i + 1);
        @(posedge clk);
        if(RD1ref !== RD1) begin 
            $display("\n\nincorrect data %h at address %h, correct data %h\n", RD1, a1, RD1ref);
            $stop();
            err_count = err_count + 1;
        end
        if(RD2ref !== RD2) begin 
            $display("\n\nincorrect data %h at address %h, correct data %h\n", RD2, a2, RD2ref);
            $stop();
            err_count = err_count + 1;
        end
      end
      if( !err_count )  $display("\n rf_riscv SUCCESS!!!\n");
      $finish();
    end
endmodule


(* STRUCTURAL_NETLIST = "yes" *)
module register_file_ref
   (clk,
    A1,
    A2,
    A3,
    WD,
    WE,
    RD1,
    RD2);
  input clk;
  input [4:0]A1;
  input [4:0]A2;
  input [4:0]A3;
  input [31:0]WD;
  input WE;
  output [31:0]RD1;
  output [31:0]RD2;

  wire \<const0> ;
  wire [4:0]A1;
  wire [4:0]A1_IBUF;
  wire [4:0]A2;
  wire [4:0]A2_IBUF;
  wire [4:0]A3;
  wire [4:0]A3_IBUF;
  wire [31:0]RD1;
  wire [31:0]RD1_OBUF;
  wire \RD1_OBUF[0]_inst_i_10_n_0 ;
  wire \RD1_OBUF[0]_inst_i_11_n_0 ;
  wire \RD1_OBUF[0]_inst_i_12_n_0 ;
  wire \RD1_OBUF[0]_inst_i_13_n_0 ;
  wire \RD1_OBUF[0]_inst_i_2_n_0 ;
  wire \RD1_OBUF[0]_inst_i_3_n_0 ;
  wire \RD1_OBUF[0]_inst_i_4_n_0 ;
  wire \RD1_OBUF[0]_inst_i_5_n_0 ;
  wire \RD1_OBUF[0]_inst_i_6_n_0 ;
  wire \RD1_OBUF[0]_inst_i_7_n_0 ;
  wire \RD1_OBUF[0]_inst_i_8_n_0 ;
  wire \RD1_OBUF[0]_inst_i_9_n_0 ;
  wire \RD1_OBUF[10]_inst_i_10_n_0 ;
  wire \RD1_OBUF[10]_inst_i_11_n_0 ;
  wire \RD1_OBUF[10]_inst_i_12_n_0 ;
  wire \RD1_OBUF[10]_inst_i_13_n_0 ;
  wire \RD1_OBUF[10]_inst_i_2_n_0 ;
  wire \RD1_OBUF[10]_inst_i_3_n_0 ;
  wire \RD1_OBUF[10]_inst_i_4_n_0 ;
  wire \RD1_OBUF[10]_inst_i_5_n_0 ;
  wire \RD1_OBUF[10]_inst_i_6_n_0 ;
  wire \RD1_OBUF[10]_inst_i_7_n_0 ;
  wire \RD1_OBUF[10]_inst_i_8_n_0 ;
  wire \RD1_OBUF[10]_inst_i_9_n_0 ;
  wire \RD1_OBUF[11]_inst_i_10_n_0 ;
  wire \RD1_OBUF[11]_inst_i_11_n_0 ;
  wire \RD1_OBUF[11]_inst_i_12_n_0 ;
  wire \RD1_OBUF[11]_inst_i_13_n_0 ;
  wire \RD1_OBUF[11]_inst_i_2_n_0 ;
  wire \RD1_OBUF[11]_inst_i_3_n_0 ;
  wire \RD1_OBUF[11]_inst_i_4_n_0 ;
  wire \RD1_OBUF[11]_inst_i_5_n_0 ;
  wire \RD1_OBUF[11]_inst_i_6_n_0 ;
  wire \RD1_OBUF[11]_inst_i_7_n_0 ;
  wire \RD1_OBUF[11]_inst_i_8_n_0 ;
  wire \RD1_OBUF[11]_inst_i_9_n_0 ;
  wire \RD1_OBUF[12]_inst_i_10_n_0 ;
  wire \RD1_OBUF[12]_inst_i_11_n_0 ;
  wire \RD1_OBUF[12]_inst_i_12_n_0 ;
  wire \RD1_OBUF[12]_inst_i_13_n_0 ;
  wire \RD1_OBUF[12]_inst_i_2_n_0 ;
  wire \RD1_OBUF[12]_inst_i_3_n_0 ;
  wire \RD1_OBUF[12]_inst_i_4_n_0 ;
  wire \RD1_OBUF[12]_inst_i_5_n_0 ;
  wire \RD1_OBUF[12]_inst_i_6_n_0 ;
  wire \RD1_OBUF[12]_inst_i_7_n_0 ;
  wire \RD1_OBUF[12]_inst_i_8_n_0 ;
  wire \RD1_OBUF[12]_inst_i_9_n_0 ;
  wire \RD1_OBUF[13]_inst_i_10_n_0 ;
  wire \RD1_OBUF[13]_inst_i_11_n_0 ;
  wire \RD1_OBUF[13]_inst_i_12_n_0 ;
  wire \RD1_OBUF[13]_inst_i_13_n_0 ;
  wire \RD1_OBUF[13]_inst_i_2_n_0 ;
  wire \RD1_OBUF[13]_inst_i_3_n_0 ;
  wire \RD1_OBUF[13]_inst_i_4_n_0 ;
  wire \RD1_OBUF[13]_inst_i_5_n_0 ;
  wire \RD1_OBUF[13]_inst_i_6_n_0 ;
  wire \RD1_OBUF[13]_inst_i_7_n_0 ;
  wire \RD1_OBUF[13]_inst_i_8_n_0 ;
  wire \RD1_OBUF[13]_inst_i_9_n_0 ;
  wire \RD1_OBUF[14]_inst_i_10_n_0 ;
  wire \RD1_OBUF[14]_inst_i_11_n_0 ;
  wire \RD1_OBUF[14]_inst_i_12_n_0 ;
  wire \RD1_OBUF[14]_inst_i_13_n_0 ;
  wire \RD1_OBUF[14]_inst_i_2_n_0 ;
  wire \RD1_OBUF[14]_inst_i_3_n_0 ;
  wire \RD1_OBUF[14]_inst_i_4_n_0 ;
  wire \RD1_OBUF[14]_inst_i_5_n_0 ;
  wire \RD1_OBUF[14]_inst_i_6_n_0 ;
  wire \RD1_OBUF[14]_inst_i_7_n_0 ;
  wire \RD1_OBUF[14]_inst_i_8_n_0 ;
  wire \RD1_OBUF[14]_inst_i_9_n_0 ;
  wire \RD1_OBUF[15]_inst_i_10_n_0 ;
  wire \RD1_OBUF[15]_inst_i_11_n_0 ;
  wire \RD1_OBUF[15]_inst_i_12_n_0 ;
  wire \RD1_OBUF[15]_inst_i_13_n_0 ;
  wire \RD1_OBUF[15]_inst_i_2_n_0 ;
  wire \RD1_OBUF[15]_inst_i_3_n_0 ;
  wire \RD1_OBUF[15]_inst_i_4_n_0 ;
  wire \RD1_OBUF[15]_inst_i_5_n_0 ;
  wire \RD1_OBUF[15]_inst_i_6_n_0 ;
  wire \RD1_OBUF[15]_inst_i_7_n_0 ;
  wire \RD1_OBUF[15]_inst_i_8_n_0 ;
  wire \RD1_OBUF[15]_inst_i_9_n_0 ;
  wire \RD1_OBUF[16]_inst_i_10_n_0 ;
  wire \RD1_OBUF[16]_inst_i_11_n_0 ;
  wire \RD1_OBUF[16]_inst_i_12_n_0 ;
  wire \RD1_OBUF[16]_inst_i_13_n_0 ;
  wire \RD1_OBUF[16]_inst_i_2_n_0 ;
  wire \RD1_OBUF[16]_inst_i_3_n_0 ;
  wire \RD1_OBUF[16]_inst_i_4_n_0 ;
  wire \RD1_OBUF[16]_inst_i_5_n_0 ;
  wire \RD1_OBUF[16]_inst_i_6_n_0 ;
  wire \RD1_OBUF[16]_inst_i_7_n_0 ;
  wire \RD1_OBUF[16]_inst_i_8_n_0 ;
  wire \RD1_OBUF[16]_inst_i_9_n_0 ;
  wire \RD1_OBUF[17]_inst_i_10_n_0 ;
  wire \RD1_OBUF[17]_inst_i_11_n_0 ;
  wire \RD1_OBUF[17]_inst_i_12_n_0 ;
  wire \RD1_OBUF[17]_inst_i_13_n_0 ;
  wire \RD1_OBUF[17]_inst_i_2_n_0 ;
  wire \RD1_OBUF[17]_inst_i_3_n_0 ;
  wire \RD1_OBUF[17]_inst_i_4_n_0 ;
  wire \RD1_OBUF[17]_inst_i_5_n_0 ;
  wire \RD1_OBUF[17]_inst_i_6_n_0 ;
  wire \RD1_OBUF[17]_inst_i_7_n_0 ;
  wire \RD1_OBUF[17]_inst_i_8_n_0 ;
  wire \RD1_OBUF[17]_inst_i_9_n_0 ;
  wire \RD1_OBUF[18]_inst_i_10_n_0 ;
  wire \RD1_OBUF[18]_inst_i_11_n_0 ;
  wire \RD1_OBUF[18]_inst_i_12_n_0 ;
  wire \RD1_OBUF[18]_inst_i_13_n_0 ;
  wire \RD1_OBUF[18]_inst_i_2_n_0 ;
  wire \RD1_OBUF[18]_inst_i_3_n_0 ;
  wire \RD1_OBUF[18]_inst_i_4_n_0 ;
  wire \RD1_OBUF[18]_inst_i_5_n_0 ;
  wire \RD1_OBUF[18]_inst_i_6_n_0 ;
  wire \RD1_OBUF[18]_inst_i_7_n_0 ;
  wire \RD1_OBUF[18]_inst_i_8_n_0 ;
  wire \RD1_OBUF[18]_inst_i_9_n_0 ;
  wire \RD1_OBUF[19]_inst_i_10_n_0 ;
  wire \RD1_OBUF[19]_inst_i_11_n_0 ;
  wire \RD1_OBUF[19]_inst_i_12_n_0 ;
  wire \RD1_OBUF[19]_inst_i_13_n_0 ;
  wire \RD1_OBUF[19]_inst_i_2_n_0 ;
  wire \RD1_OBUF[19]_inst_i_3_n_0 ;
  wire \RD1_OBUF[19]_inst_i_4_n_0 ;
  wire \RD1_OBUF[19]_inst_i_5_n_0 ;
  wire \RD1_OBUF[19]_inst_i_6_n_0 ;
  wire \RD1_OBUF[19]_inst_i_7_n_0 ;
  wire \RD1_OBUF[19]_inst_i_8_n_0 ;
  wire \RD1_OBUF[19]_inst_i_9_n_0 ;
  wire \RD1_OBUF[1]_inst_i_10_n_0 ;
  wire \RD1_OBUF[1]_inst_i_11_n_0 ;
  wire \RD1_OBUF[1]_inst_i_12_n_0 ;
  wire \RD1_OBUF[1]_inst_i_13_n_0 ;
  wire \RD1_OBUF[1]_inst_i_2_n_0 ;
  wire \RD1_OBUF[1]_inst_i_3_n_0 ;
  wire \RD1_OBUF[1]_inst_i_4_n_0 ;
  wire \RD1_OBUF[1]_inst_i_5_n_0 ;
  wire \RD1_OBUF[1]_inst_i_6_n_0 ;
  wire \RD1_OBUF[1]_inst_i_7_n_0 ;
  wire \RD1_OBUF[1]_inst_i_8_n_0 ;
  wire \RD1_OBUF[1]_inst_i_9_n_0 ;
  wire \RD1_OBUF[20]_inst_i_10_n_0 ;
  wire \RD1_OBUF[20]_inst_i_11_n_0 ;
  wire \RD1_OBUF[20]_inst_i_12_n_0 ;
  wire \RD1_OBUF[20]_inst_i_13_n_0 ;
  wire \RD1_OBUF[20]_inst_i_2_n_0 ;
  wire \RD1_OBUF[20]_inst_i_3_n_0 ;
  wire \RD1_OBUF[20]_inst_i_4_n_0 ;
  wire \RD1_OBUF[20]_inst_i_5_n_0 ;
  wire \RD1_OBUF[20]_inst_i_6_n_0 ;
  wire \RD1_OBUF[20]_inst_i_7_n_0 ;
  wire \RD1_OBUF[20]_inst_i_8_n_0 ;
  wire \RD1_OBUF[20]_inst_i_9_n_0 ;
  wire \RD1_OBUF[21]_inst_i_10_n_0 ;
  wire \RD1_OBUF[21]_inst_i_11_n_0 ;
  wire \RD1_OBUF[21]_inst_i_12_n_0 ;
  wire \RD1_OBUF[21]_inst_i_13_n_0 ;
  wire \RD1_OBUF[21]_inst_i_2_n_0 ;
  wire \RD1_OBUF[21]_inst_i_3_n_0 ;
  wire \RD1_OBUF[21]_inst_i_4_n_0 ;
  wire \RD1_OBUF[21]_inst_i_5_n_0 ;
  wire \RD1_OBUF[21]_inst_i_6_n_0 ;
  wire \RD1_OBUF[21]_inst_i_7_n_0 ;
  wire \RD1_OBUF[21]_inst_i_8_n_0 ;
  wire \RD1_OBUF[21]_inst_i_9_n_0 ;
  wire \RD1_OBUF[22]_inst_i_10_n_0 ;
  wire \RD1_OBUF[22]_inst_i_11_n_0 ;
  wire \RD1_OBUF[22]_inst_i_12_n_0 ;
  wire \RD1_OBUF[22]_inst_i_13_n_0 ;
  wire \RD1_OBUF[22]_inst_i_2_n_0 ;
  wire \RD1_OBUF[22]_inst_i_3_n_0 ;
  wire \RD1_OBUF[22]_inst_i_4_n_0 ;
  wire \RD1_OBUF[22]_inst_i_5_n_0 ;
  wire \RD1_OBUF[22]_inst_i_6_n_0 ;
  wire \RD1_OBUF[22]_inst_i_7_n_0 ;
  wire \RD1_OBUF[22]_inst_i_8_n_0 ;
  wire \RD1_OBUF[22]_inst_i_9_n_0 ;
  wire \RD1_OBUF[23]_inst_i_10_n_0 ;
  wire \RD1_OBUF[23]_inst_i_11_n_0 ;
  wire \RD1_OBUF[23]_inst_i_12_n_0 ;
  wire \RD1_OBUF[23]_inst_i_13_n_0 ;
  wire \RD1_OBUF[23]_inst_i_2_n_0 ;
  wire \RD1_OBUF[23]_inst_i_3_n_0 ;
  wire \RD1_OBUF[23]_inst_i_4_n_0 ;
  wire \RD1_OBUF[23]_inst_i_5_n_0 ;
  wire \RD1_OBUF[23]_inst_i_6_n_0 ;
  wire \RD1_OBUF[23]_inst_i_7_n_0 ;
  wire \RD1_OBUF[23]_inst_i_8_n_0 ;
  wire \RD1_OBUF[23]_inst_i_9_n_0 ;
  wire \RD1_OBUF[24]_inst_i_10_n_0 ;
  wire \RD1_OBUF[24]_inst_i_11_n_0 ;
  wire \RD1_OBUF[24]_inst_i_12_n_0 ;
  wire \RD1_OBUF[24]_inst_i_13_n_0 ;
  wire \RD1_OBUF[24]_inst_i_2_n_0 ;
  wire \RD1_OBUF[24]_inst_i_3_n_0 ;
  wire \RD1_OBUF[24]_inst_i_4_n_0 ;
  wire \RD1_OBUF[24]_inst_i_5_n_0 ;
  wire \RD1_OBUF[24]_inst_i_6_n_0 ;
  wire \RD1_OBUF[24]_inst_i_7_n_0 ;
  wire \RD1_OBUF[24]_inst_i_8_n_0 ;
  wire \RD1_OBUF[24]_inst_i_9_n_0 ;
  wire \RD1_OBUF[25]_inst_i_10_n_0 ;
  wire \RD1_OBUF[25]_inst_i_11_n_0 ;
  wire \RD1_OBUF[25]_inst_i_12_n_0 ;
  wire \RD1_OBUF[25]_inst_i_13_n_0 ;
  wire \RD1_OBUF[25]_inst_i_2_n_0 ;
  wire \RD1_OBUF[25]_inst_i_3_n_0 ;
  wire \RD1_OBUF[25]_inst_i_4_n_0 ;
  wire \RD1_OBUF[25]_inst_i_5_n_0 ;
  wire \RD1_OBUF[25]_inst_i_6_n_0 ;
  wire \RD1_OBUF[25]_inst_i_7_n_0 ;
  wire \RD1_OBUF[25]_inst_i_8_n_0 ;
  wire \RD1_OBUF[25]_inst_i_9_n_0 ;
  wire \RD1_OBUF[26]_inst_i_10_n_0 ;
  wire \RD1_OBUF[26]_inst_i_11_n_0 ;
  wire \RD1_OBUF[26]_inst_i_12_n_0 ;
  wire \RD1_OBUF[26]_inst_i_13_n_0 ;
  wire \RD1_OBUF[26]_inst_i_2_n_0 ;
  wire \RD1_OBUF[26]_inst_i_3_n_0 ;
  wire \RD1_OBUF[26]_inst_i_4_n_0 ;
  wire \RD1_OBUF[26]_inst_i_5_n_0 ;
  wire \RD1_OBUF[26]_inst_i_6_n_0 ;
  wire \RD1_OBUF[26]_inst_i_7_n_0 ;
  wire \RD1_OBUF[26]_inst_i_8_n_0 ;
  wire \RD1_OBUF[26]_inst_i_9_n_0 ;
  wire \RD1_OBUF[27]_inst_i_10_n_0 ;
  wire \RD1_OBUF[27]_inst_i_11_n_0 ;
  wire \RD1_OBUF[27]_inst_i_12_n_0 ;
  wire \RD1_OBUF[27]_inst_i_13_n_0 ;
  wire \RD1_OBUF[27]_inst_i_2_n_0 ;
  wire \RD1_OBUF[27]_inst_i_3_n_0 ;
  wire \RD1_OBUF[27]_inst_i_4_n_0 ;
  wire \RD1_OBUF[27]_inst_i_5_n_0 ;
  wire \RD1_OBUF[27]_inst_i_6_n_0 ;
  wire \RD1_OBUF[27]_inst_i_7_n_0 ;
  wire \RD1_OBUF[27]_inst_i_8_n_0 ;
  wire \RD1_OBUF[27]_inst_i_9_n_0 ;
  wire \RD1_OBUF[28]_inst_i_10_n_0 ;
  wire \RD1_OBUF[28]_inst_i_11_n_0 ;
  wire \RD1_OBUF[28]_inst_i_12_n_0 ;
  wire \RD1_OBUF[28]_inst_i_13_n_0 ;
  wire \RD1_OBUF[28]_inst_i_2_n_0 ;
  wire \RD1_OBUF[28]_inst_i_3_n_0 ;
  wire \RD1_OBUF[28]_inst_i_4_n_0 ;
  wire \RD1_OBUF[28]_inst_i_5_n_0 ;
  wire \RD1_OBUF[28]_inst_i_6_n_0 ;
  wire \RD1_OBUF[28]_inst_i_7_n_0 ;
  wire \RD1_OBUF[28]_inst_i_8_n_0 ;
  wire \RD1_OBUF[28]_inst_i_9_n_0 ;
  wire \RD1_OBUF[29]_inst_i_10_n_0 ;
  wire \RD1_OBUF[29]_inst_i_11_n_0 ;
  wire \RD1_OBUF[29]_inst_i_12_n_0 ;
  wire \RD1_OBUF[29]_inst_i_13_n_0 ;
  wire \RD1_OBUF[29]_inst_i_2_n_0 ;
  wire \RD1_OBUF[29]_inst_i_3_n_0 ;
  wire \RD1_OBUF[29]_inst_i_4_n_0 ;
  wire \RD1_OBUF[29]_inst_i_5_n_0 ;
  wire \RD1_OBUF[29]_inst_i_6_n_0 ;
  wire \RD1_OBUF[29]_inst_i_7_n_0 ;
  wire \RD1_OBUF[29]_inst_i_8_n_0 ;
  wire \RD1_OBUF[29]_inst_i_9_n_0 ;
  wire \RD1_OBUF[2]_inst_i_10_n_0 ;
  wire \RD1_OBUF[2]_inst_i_11_n_0 ;
  wire \RD1_OBUF[2]_inst_i_12_n_0 ;
  wire \RD1_OBUF[2]_inst_i_13_n_0 ;
  wire \RD1_OBUF[2]_inst_i_2_n_0 ;
  wire \RD1_OBUF[2]_inst_i_3_n_0 ;
  wire \RD1_OBUF[2]_inst_i_4_n_0 ;
  wire \RD1_OBUF[2]_inst_i_5_n_0 ;
  wire \RD1_OBUF[2]_inst_i_6_n_0 ;
  wire \RD1_OBUF[2]_inst_i_7_n_0 ;
  wire \RD1_OBUF[2]_inst_i_8_n_0 ;
  wire \RD1_OBUF[2]_inst_i_9_n_0 ;
  wire \RD1_OBUF[30]_inst_i_10_n_0 ;
  wire \RD1_OBUF[30]_inst_i_11_n_0 ;
  wire \RD1_OBUF[30]_inst_i_12_n_0 ;
  wire \RD1_OBUF[30]_inst_i_13_n_0 ;
  wire \RD1_OBUF[30]_inst_i_2_n_0 ;
  wire \RD1_OBUF[30]_inst_i_3_n_0 ;
  wire \RD1_OBUF[30]_inst_i_4_n_0 ;
  wire \RD1_OBUF[30]_inst_i_5_n_0 ;
  wire \RD1_OBUF[30]_inst_i_6_n_0 ;
  wire \RD1_OBUF[30]_inst_i_7_n_0 ;
  wire \RD1_OBUF[30]_inst_i_8_n_0 ;
  wire \RD1_OBUF[30]_inst_i_9_n_0 ;
  wire \RD1_OBUF[31]_inst_i_10_n_0 ;
  wire \RD1_OBUF[31]_inst_i_11_n_0 ;
  wire \RD1_OBUF[31]_inst_i_12_n_0 ;
  wire \RD1_OBUF[31]_inst_i_13_n_0 ;
  wire \RD1_OBUF[31]_inst_i_2_n_0 ;
  wire \RD1_OBUF[31]_inst_i_3_n_0 ;
  wire \RD1_OBUF[31]_inst_i_4_n_0 ;
  wire \RD1_OBUF[31]_inst_i_5_n_0 ;
  wire \RD1_OBUF[31]_inst_i_6_n_0 ;
  wire \RD1_OBUF[31]_inst_i_7_n_0 ;
  wire \RD1_OBUF[31]_inst_i_8_n_0 ;
  wire \RD1_OBUF[31]_inst_i_9_n_0 ;
  wire \RD1_OBUF[3]_inst_i_10_n_0 ;
  wire \RD1_OBUF[3]_inst_i_11_n_0 ;
  wire \RD1_OBUF[3]_inst_i_12_n_0 ;
  wire \RD1_OBUF[3]_inst_i_13_n_0 ;
  wire \RD1_OBUF[3]_inst_i_2_n_0 ;
  wire \RD1_OBUF[3]_inst_i_3_n_0 ;
  wire \RD1_OBUF[3]_inst_i_4_n_0 ;
  wire \RD1_OBUF[3]_inst_i_5_n_0 ;
  wire \RD1_OBUF[3]_inst_i_6_n_0 ;
  wire \RD1_OBUF[3]_inst_i_7_n_0 ;
  wire \RD1_OBUF[3]_inst_i_8_n_0 ;
  wire \RD1_OBUF[3]_inst_i_9_n_0 ;
  wire \RD1_OBUF[4]_inst_i_10_n_0 ;
  wire \RD1_OBUF[4]_inst_i_11_n_0 ;
  wire \RD1_OBUF[4]_inst_i_12_n_0 ;
  wire \RD1_OBUF[4]_inst_i_13_n_0 ;
  wire \RD1_OBUF[4]_inst_i_2_n_0 ;
  wire \RD1_OBUF[4]_inst_i_3_n_0 ;
  wire \RD1_OBUF[4]_inst_i_4_n_0 ;
  wire \RD1_OBUF[4]_inst_i_5_n_0 ;
  wire \RD1_OBUF[4]_inst_i_6_n_0 ;
  wire \RD1_OBUF[4]_inst_i_7_n_0 ;
  wire \RD1_OBUF[4]_inst_i_8_n_0 ;
  wire \RD1_OBUF[4]_inst_i_9_n_0 ;
  wire \RD1_OBUF[5]_inst_i_10_n_0 ;
  wire \RD1_OBUF[5]_inst_i_11_n_0 ;
  wire \RD1_OBUF[5]_inst_i_12_n_0 ;
  wire \RD1_OBUF[5]_inst_i_13_n_0 ;
  wire \RD1_OBUF[5]_inst_i_2_n_0 ;
  wire \RD1_OBUF[5]_inst_i_3_n_0 ;
  wire \RD1_OBUF[5]_inst_i_4_n_0 ;
  wire \RD1_OBUF[5]_inst_i_5_n_0 ;
  wire \RD1_OBUF[5]_inst_i_6_n_0 ;
  wire \RD1_OBUF[5]_inst_i_7_n_0 ;
  wire \RD1_OBUF[5]_inst_i_8_n_0 ;
  wire \RD1_OBUF[5]_inst_i_9_n_0 ;
  wire \RD1_OBUF[6]_inst_i_10_n_0 ;
  wire \RD1_OBUF[6]_inst_i_11_n_0 ;
  wire \RD1_OBUF[6]_inst_i_12_n_0 ;
  wire \RD1_OBUF[6]_inst_i_13_n_0 ;
  wire \RD1_OBUF[6]_inst_i_2_n_0 ;
  wire \RD1_OBUF[6]_inst_i_3_n_0 ;
  wire \RD1_OBUF[6]_inst_i_4_n_0 ;
  wire \RD1_OBUF[6]_inst_i_5_n_0 ;
  wire \RD1_OBUF[6]_inst_i_6_n_0 ;
  wire \RD1_OBUF[6]_inst_i_7_n_0 ;
  wire \RD1_OBUF[6]_inst_i_8_n_0 ;
  wire \RD1_OBUF[6]_inst_i_9_n_0 ;
  wire \RD1_OBUF[7]_inst_i_10_n_0 ;
  wire \RD1_OBUF[7]_inst_i_11_n_0 ;
  wire \RD1_OBUF[7]_inst_i_12_n_0 ;
  wire \RD1_OBUF[7]_inst_i_13_n_0 ;
  wire \RD1_OBUF[7]_inst_i_2_n_0 ;
  wire \RD1_OBUF[7]_inst_i_3_n_0 ;
  wire \RD1_OBUF[7]_inst_i_4_n_0 ;
  wire \RD1_OBUF[7]_inst_i_5_n_0 ;
  wire \RD1_OBUF[7]_inst_i_6_n_0 ;
  wire \RD1_OBUF[7]_inst_i_7_n_0 ;
  wire \RD1_OBUF[7]_inst_i_8_n_0 ;
  wire \RD1_OBUF[7]_inst_i_9_n_0 ;
  wire \RD1_OBUF[8]_inst_i_10_n_0 ;
  wire \RD1_OBUF[8]_inst_i_11_n_0 ;
  wire \RD1_OBUF[8]_inst_i_12_n_0 ;
  wire \RD1_OBUF[8]_inst_i_13_n_0 ;
  wire \RD1_OBUF[8]_inst_i_2_n_0 ;
  wire \RD1_OBUF[8]_inst_i_3_n_0 ;
  wire \RD1_OBUF[8]_inst_i_4_n_0 ;
  wire \RD1_OBUF[8]_inst_i_5_n_0 ;
  wire \RD1_OBUF[8]_inst_i_6_n_0 ;
  wire \RD1_OBUF[8]_inst_i_7_n_0 ;
  wire \RD1_OBUF[8]_inst_i_8_n_0 ;
  wire \RD1_OBUF[8]_inst_i_9_n_0 ;
  wire \RD1_OBUF[9]_inst_i_10_n_0 ;
  wire \RD1_OBUF[9]_inst_i_11_n_0 ;
  wire \RD1_OBUF[9]_inst_i_12_n_0 ;
  wire \RD1_OBUF[9]_inst_i_13_n_0 ;
  wire \RD1_OBUF[9]_inst_i_2_n_0 ;
  wire \RD1_OBUF[9]_inst_i_3_n_0 ;
  wire \RD1_OBUF[9]_inst_i_4_n_0 ;
  wire \RD1_OBUF[9]_inst_i_5_n_0 ;
  wire \RD1_OBUF[9]_inst_i_6_n_0 ;
  wire \RD1_OBUF[9]_inst_i_7_n_0 ;
  wire \RD1_OBUF[9]_inst_i_8_n_0 ;
  wire \RD1_OBUF[9]_inst_i_9_n_0 ;
  wire [31:0]RD2;
  wire [31:0]RD2_OBUF;
  wire \RD2_OBUF[0]_inst_i_10_n_0 ;
  wire \RD2_OBUF[0]_inst_i_11_n_0 ;
  wire \RD2_OBUF[0]_inst_i_12_n_0 ;
  wire \RD2_OBUF[0]_inst_i_13_n_0 ;
  wire \RD2_OBUF[0]_inst_i_2_n_0 ;
  wire \RD2_OBUF[0]_inst_i_3_n_0 ;
  wire \RD2_OBUF[0]_inst_i_4_n_0 ;
  wire \RD2_OBUF[0]_inst_i_5_n_0 ;
  wire \RD2_OBUF[0]_inst_i_6_n_0 ;
  wire \RD2_OBUF[0]_inst_i_7_n_0 ;
  wire \RD2_OBUF[0]_inst_i_8_n_0 ;
  wire \RD2_OBUF[0]_inst_i_9_n_0 ;
  wire \RD2_OBUF[10]_inst_i_10_n_0 ;
  wire \RD2_OBUF[10]_inst_i_11_n_0 ;
  wire \RD2_OBUF[10]_inst_i_12_n_0 ;
  wire \RD2_OBUF[10]_inst_i_13_n_0 ;
  wire \RD2_OBUF[10]_inst_i_2_n_0 ;
  wire \RD2_OBUF[10]_inst_i_3_n_0 ;
  wire \RD2_OBUF[10]_inst_i_4_n_0 ;
  wire \RD2_OBUF[10]_inst_i_5_n_0 ;
  wire \RD2_OBUF[10]_inst_i_6_n_0 ;
  wire \RD2_OBUF[10]_inst_i_7_n_0 ;
  wire \RD2_OBUF[10]_inst_i_8_n_0 ;
  wire \RD2_OBUF[10]_inst_i_9_n_0 ;
  wire \RD2_OBUF[11]_inst_i_10_n_0 ;
  wire \RD2_OBUF[11]_inst_i_11_n_0 ;
  wire \RD2_OBUF[11]_inst_i_12_n_0 ;
  wire \RD2_OBUF[11]_inst_i_13_n_0 ;
  wire \RD2_OBUF[11]_inst_i_2_n_0 ;
  wire \RD2_OBUF[11]_inst_i_3_n_0 ;
  wire \RD2_OBUF[11]_inst_i_4_n_0 ;
  wire \RD2_OBUF[11]_inst_i_5_n_0 ;
  wire \RD2_OBUF[11]_inst_i_6_n_0 ;
  wire \RD2_OBUF[11]_inst_i_7_n_0 ;
  wire \RD2_OBUF[11]_inst_i_8_n_0 ;
  wire \RD2_OBUF[11]_inst_i_9_n_0 ;
  wire \RD2_OBUF[12]_inst_i_10_n_0 ;
  wire \RD2_OBUF[12]_inst_i_11_n_0 ;
  wire \RD2_OBUF[12]_inst_i_12_n_0 ;
  wire \RD2_OBUF[12]_inst_i_13_n_0 ;
  wire \RD2_OBUF[12]_inst_i_2_n_0 ;
  wire \RD2_OBUF[12]_inst_i_3_n_0 ;
  wire \RD2_OBUF[12]_inst_i_4_n_0 ;
  wire \RD2_OBUF[12]_inst_i_5_n_0 ;
  wire \RD2_OBUF[12]_inst_i_6_n_0 ;
  wire \RD2_OBUF[12]_inst_i_7_n_0 ;
  wire \RD2_OBUF[12]_inst_i_8_n_0 ;
  wire \RD2_OBUF[12]_inst_i_9_n_0 ;
  wire \RD2_OBUF[13]_inst_i_10_n_0 ;
  wire \RD2_OBUF[13]_inst_i_11_n_0 ;
  wire \RD2_OBUF[13]_inst_i_12_n_0 ;
  wire \RD2_OBUF[13]_inst_i_13_n_0 ;
  wire \RD2_OBUF[13]_inst_i_2_n_0 ;
  wire \RD2_OBUF[13]_inst_i_3_n_0 ;
  wire \RD2_OBUF[13]_inst_i_4_n_0 ;
  wire \RD2_OBUF[13]_inst_i_5_n_0 ;
  wire \RD2_OBUF[13]_inst_i_6_n_0 ;
  wire \RD2_OBUF[13]_inst_i_7_n_0 ;
  wire \RD2_OBUF[13]_inst_i_8_n_0 ;
  wire \RD2_OBUF[13]_inst_i_9_n_0 ;
  wire \RD2_OBUF[14]_inst_i_10_n_0 ;
  wire \RD2_OBUF[14]_inst_i_11_n_0 ;
  wire \RD2_OBUF[14]_inst_i_12_n_0 ;
  wire \RD2_OBUF[14]_inst_i_13_n_0 ;
  wire \RD2_OBUF[14]_inst_i_2_n_0 ;
  wire \RD2_OBUF[14]_inst_i_3_n_0 ;
  wire \RD2_OBUF[14]_inst_i_4_n_0 ;
  wire \RD2_OBUF[14]_inst_i_5_n_0 ;
  wire \RD2_OBUF[14]_inst_i_6_n_0 ;
  wire \RD2_OBUF[14]_inst_i_7_n_0 ;
  wire \RD2_OBUF[14]_inst_i_8_n_0 ;
  wire \RD2_OBUF[14]_inst_i_9_n_0 ;
  wire \RD2_OBUF[15]_inst_i_10_n_0 ;
  wire \RD2_OBUF[15]_inst_i_11_n_0 ;
  wire \RD2_OBUF[15]_inst_i_12_n_0 ;
  wire \RD2_OBUF[15]_inst_i_13_n_0 ;
  wire \RD2_OBUF[15]_inst_i_2_n_0 ;
  wire \RD2_OBUF[15]_inst_i_3_n_0 ;
  wire \RD2_OBUF[15]_inst_i_4_n_0 ;
  wire \RD2_OBUF[15]_inst_i_5_n_0 ;
  wire \RD2_OBUF[15]_inst_i_6_n_0 ;
  wire \RD2_OBUF[15]_inst_i_7_n_0 ;
  wire \RD2_OBUF[15]_inst_i_8_n_0 ;
  wire \RD2_OBUF[15]_inst_i_9_n_0 ;
  wire \RD2_OBUF[16]_inst_i_10_n_0 ;
  wire \RD2_OBUF[16]_inst_i_11_n_0 ;
  wire \RD2_OBUF[16]_inst_i_12_n_0 ;
  wire \RD2_OBUF[16]_inst_i_13_n_0 ;
  wire \RD2_OBUF[16]_inst_i_2_n_0 ;
  wire \RD2_OBUF[16]_inst_i_3_n_0 ;
  wire \RD2_OBUF[16]_inst_i_4_n_0 ;
  wire \RD2_OBUF[16]_inst_i_5_n_0 ;
  wire \RD2_OBUF[16]_inst_i_6_n_0 ;
  wire \RD2_OBUF[16]_inst_i_7_n_0 ;
  wire \RD2_OBUF[16]_inst_i_8_n_0 ;
  wire \RD2_OBUF[16]_inst_i_9_n_0 ;
  wire \RD2_OBUF[17]_inst_i_10_n_0 ;
  wire \RD2_OBUF[17]_inst_i_11_n_0 ;
  wire \RD2_OBUF[17]_inst_i_12_n_0 ;
  wire \RD2_OBUF[17]_inst_i_13_n_0 ;
  wire \RD2_OBUF[17]_inst_i_2_n_0 ;
  wire \RD2_OBUF[17]_inst_i_3_n_0 ;
  wire \RD2_OBUF[17]_inst_i_4_n_0 ;
  wire \RD2_OBUF[17]_inst_i_5_n_0 ;
  wire \RD2_OBUF[17]_inst_i_6_n_0 ;
  wire \RD2_OBUF[17]_inst_i_7_n_0 ;
  wire \RD2_OBUF[17]_inst_i_8_n_0 ;
  wire \RD2_OBUF[17]_inst_i_9_n_0 ;
  wire \RD2_OBUF[18]_inst_i_10_n_0 ;
  wire \RD2_OBUF[18]_inst_i_11_n_0 ;
  wire \RD2_OBUF[18]_inst_i_12_n_0 ;
  wire \RD2_OBUF[18]_inst_i_13_n_0 ;
  wire \RD2_OBUF[18]_inst_i_2_n_0 ;
  wire \RD2_OBUF[18]_inst_i_3_n_0 ;
  wire \RD2_OBUF[18]_inst_i_4_n_0 ;
  wire \RD2_OBUF[18]_inst_i_5_n_0 ;
  wire \RD2_OBUF[18]_inst_i_6_n_0 ;
  wire \RD2_OBUF[18]_inst_i_7_n_0 ;
  wire \RD2_OBUF[18]_inst_i_8_n_0 ;
  wire \RD2_OBUF[18]_inst_i_9_n_0 ;
  wire \RD2_OBUF[19]_inst_i_10_n_0 ;
  wire \RD2_OBUF[19]_inst_i_11_n_0 ;
  wire \RD2_OBUF[19]_inst_i_12_n_0 ;
  wire \RD2_OBUF[19]_inst_i_13_n_0 ;
  wire \RD2_OBUF[19]_inst_i_2_n_0 ;
  wire \RD2_OBUF[19]_inst_i_3_n_0 ;
  wire \RD2_OBUF[19]_inst_i_4_n_0 ;
  wire \RD2_OBUF[19]_inst_i_5_n_0 ;
  wire \RD2_OBUF[19]_inst_i_6_n_0 ;
  wire \RD2_OBUF[19]_inst_i_7_n_0 ;
  wire \RD2_OBUF[19]_inst_i_8_n_0 ;
  wire \RD2_OBUF[19]_inst_i_9_n_0 ;
  wire \RD2_OBUF[1]_inst_i_10_n_0 ;
  wire \RD2_OBUF[1]_inst_i_11_n_0 ;
  wire \RD2_OBUF[1]_inst_i_12_n_0 ;
  wire \RD2_OBUF[1]_inst_i_13_n_0 ;
  wire \RD2_OBUF[1]_inst_i_2_n_0 ;
  wire \RD2_OBUF[1]_inst_i_3_n_0 ;
  wire \RD2_OBUF[1]_inst_i_4_n_0 ;
  wire \RD2_OBUF[1]_inst_i_5_n_0 ;
  wire \RD2_OBUF[1]_inst_i_6_n_0 ;
  wire \RD2_OBUF[1]_inst_i_7_n_0 ;
  wire \RD2_OBUF[1]_inst_i_8_n_0 ;
  wire \RD2_OBUF[1]_inst_i_9_n_0 ;
  wire \RD2_OBUF[20]_inst_i_10_n_0 ;
  wire \RD2_OBUF[20]_inst_i_11_n_0 ;
  wire \RD2_OBUF[20]_inst_i_12_n_0 ;
  wire \RD2_OBUF[20]_inst_i_13_n_0 ;
  wire \RD2_OBUF[20]_inst_i_2_n_0 ;
  wire \RD2_OBUF[20]_inst_i_3_n_0 ;
  wire \RD2_OBUF[20]_inst_i_4_n_0 ;
  wire \RD2_OBUF[20]_inst_i_5_n_0 ;
  wire \RD2_OBUF[20]_inst_i_6_n_0 ;
  wire \RD2_OBUF[20]_inst_i_7_n_0 ;
  wire \RD2_OBUF[20]_inst_i_8_n_0 ;
  wire \RD2_OBUF[20]_inst_i_9_n_0 ;
  wire \RD2_OBUF[21]_inst_i_10_n_0 ;
  wire \RD2_OBUF[21]_inst_i_11_n_0 ;
  wire \RD2_OBUF[21]_inst_i_12_n_0 ;
  wire \RD2_OBUF[21]_inst_i_13_n_0 ;
  wire \RD2_OBUF[21]_inst_i_2_n_0 ;
  wire \RD2_OBUF[21]_inst_i_3_n_0 ;
  wire \RD2_OBUF[21]_inst_i_4_n_0 ;
  wire \RD2_OBUF[21]_inst_i_5_n_0 ;
  wire \RD2_OBUF[21]_inst_i_6_n_0 ;
  wire \RD2_OBUF[21]_inst_i_7_n_0 ;
  wire \RD2_OBUF[21]_inst_i_8_n_0 ;
  wire \RD2_OBUF[21]_inst_i_9_n_0 ;
  wire \RD2_OBUF[22]_inst_i_10_n_0 ;
  wire \RD2_OBUF[22]_inst_i_11_n_0 ;
  wire \RD2_OBUF[22]_inst_i_12_n_0 ;
  wire \RD2_OBUF[22]_inst_i_13_n_0 ;
  wire \RD2_OBUF[22]_inst_i_2_n_0 ;
  wire \RD2_OBUF[22]_inst_i_3_n_0 ;
  wire \RD2_OBUF[22]_inst_i_4_n_0 ;
  wire \RD2_OBUF[22]_inst_i_5_n_0 ;
  wire \RD2_OBUF[22]_inst_i_6_n_0 ;
  wire \RD2_OBUF[22]_inst_i_7_n_0 ;
  wire \RD2_OBUF[22]_inst_i_8_n_0 ;
  wire \RD2_OBUF[22]_inst_i_9_n_0 ;
  wire \RD2_OBUF[23]_inst_i_10_n_0 ;
  wire \RD2_OBUF[23]_inst_i_11_n_0 ;
  wire \RD2_OBUF[23]_inst_i_12_n_0 ;
  wire \RD2_OBUF[23]_inst_i_13_n_0 ;
  wire \RD2_OBUF[23]_inst_i_2_n_0 ;
  wire \RD2_OBUF[23]_inst_i_3_n_0 ;
  wire \RD2_OBUF[23]_inst_i_4_n_0 ;
  wire \RD2_OBUF[23]_inst_i_5_n_0 ;
  wire \RD2_OBUF[23]_inst_i_6_n_0 ;
  wire \RD2_OBUF[23]_inst_i_7_n_0 ;
  wire \RD2_OBUF[23]_inst_i_8_n_0 ;
  wire \RD2_OBUF[23]_inst_i_9_n_0 ;
  wire \RD2_OBUF[24]_inst_i_10_n_0 ;
  wire \RD2_OBUF[24]_inst_i_11_n_0 ;
  wire \RD2_OBUF[24]_inst_i_12_n_0 ;
  wire \RD2_OBUF[24]_inst_i_13_n_0 ;
  wire \RD2_OBUF[24]_inst_i_2_n_0 ;
  wire \RD2_OBUF[24]_inst_i_3_n_0 ;
  wire \RD2_OBUF[24]_inst_i_4_n_0 ;
  wire \RD2_OBUF[24]_inst_i_5_n_0 ;
  wire \RD2_OBUF[24]_inst_i_6_n_0 ;
  wire \RD2_OBUF[24]_inst_i_7_n_0 ;
  wire \RD2_OBUF[24]_inst_i_8_n_0 ;
  wire \RD2_OBUF[24]_inst_i_9_n_0 ;
  wire \RD2_OBUF[25]_inst_i_10_n_0 ;
  wire \RD2_OBUF[25]_inst_i_11_n_0 ;
  wire \RD2_OBUF[25]_inst_i_12_n_0 ;
  wire \RD2_OBUF[25]_inst_i_13_n_0 ;
  wire \RD2_OBUF[25]_inst_i_2_n_0 ;
  wire \RD2_OBUF[25]_inst_i_3_n_0 ;
  wire \RD2_OBUF[25]_inst_i_4_n_0 ;
  wire \RD2_OBUF[25]_inst_i_5_n_0 ;
  wire \RD2_OBUF[25]_inst_i_6_n_0 ;
  wire \RD2_OBUF[25]_inst_i_7_n_0 ;
  wire \RD2_OBUF[25]_inst_i_8_n_0 ;
  wire \RD2_OBUF[25]_inst_i_9_n_0 ;
  wire \RD2_OBUF[26]_inst_i_10_n_0 ;
  wire \RD2_OBUF[26]_inst_i_11_n_0 ;
  wire \RD2_OBUF[26]_inst_i_12_n_0 ;
  wire \RD2_OBUF[26]_inst_i_13_n_0 ;
  wire \RD2_OBUF[26]_inst_i_2_n_0 ;
  wire \RD2_OBUF[26]_inst_i_3_n_0 ;
  wire \RD2_OBUF[26]_inst_i_4_n_0 ;
  wire \RD2_OBUF[26]_inst_i_5_n_0 ;
  wire \RD2_OBUF[26]_inst_i_6_n_0 ;
  wire \RD2_OBUF[26]_inst_i_7_n_0 ;
  wire \RD2_OBUF[26]_inst_i_8_n_0 ;
  wire \RD2_OBUF[26]_inst_i_9_n_0 ;
  wire \RD2_OBUF[27]_inst_i_10_n_0 ;
  wire \RD2_OBUF[27]_inst_i_11_n_0 ;
  wire \RD2_OBUF[27]_inst_i_12_n_0 ;
  wire \RD2_OBUF[27]_inst_i_13_n_0 ;
  wire \RD2_OBUF[27]_inst_i_2_n_0 ;
  wire \RD2_OBUF[27]_inst_i_3_n_0 ;
  wire \RD2_OBUF[27]_inst_i_4_n_0 ;
  wire \RD2_OBUF[27]_inst_i_5_n_0 ;
  wire \RD2_OBUF[27]_inst_i_6_n_0 ;
  wire \RD2_OBUF[27]_inst_i_7_n_0 ;
  wire \RD2_OBUF[27]_inst_i_8_n_0 ;
  wire \RD2_OBUF[27]_inst_i_9_n_0 ;
  wire \RD2_OBUF[28]_inst_i_10_n_0 ;
  wire \RD2_OBUF[28]_inst_i_11_n_0 ;
  wire \RD2_OBUF[28]_inst_i_12_n_0 ;
  wire \RD2_OBUF[28]_inst_i_13_n_0 ;
  wire \RD2_OBUF[28]_inst_i_2_n_0 ;
  wire \RD2_OBUF[28]_inst_i_3_n_0 ;
  wire \RD2_OBUF[28]_inst_i_4_n_0 ;
  wire \RD2_OBUF[28]_inst_i_5_n_0 ;
  wire \RD2_OBUF[28]_inst_i_6_n_0 ;
  wire \RD2_OBUF[28]_inst_i_7_n_0 ;
  wire \RD2_OBUF[28]_inst_i_8_n_0 ;
  wire \RD2_OBUF[28]_inst_i_9_n_0 ;
  wire \RD2_OBUF[29]_inst_i_10_n_0 ;
  wire \RD2_OBUF[29]_inst_i_11_n_0 ;
  wire \RD2_OBUF[29]_inst_i_12_n_0 ;
  wire \RD2_OBUF[29]_inst_i_13_n_0 ;
  wire \RD2_OBUF[29]_inst_i_2_n_0 ;
  wire \RD2_OBUF[29]_inst_i_3_n_0 ;
  wire \RD2_OBUF[29]_inst_i_4_n_0 ;
  wire \RD2_OBUF[29]_inst_i_5_n_0 ;
  wire \RD2_OBUF[29]_inst_i_6_n_0 ;
  wire \RD2_OBUF[29]_inst_i_7_n_0 ;
  wire \RD2_OBUF[29]_inst_i_8_n_0 ;
  wire \RD2_OBUF[29]_inst_i_9_n_0 ;
  wire \RD2_OBUF[2]_inst_i_10_n_0 ;
  wire \RD2_OBUF[2]_inst_i_11_n_0 ;
  wire \RD2_OBUF[2]_inst_i_12_n_0 ;
  wire \RD2_OBUF[2]_inst_i_13_n_0 ;
  wire \RD2_OBUF[2]_inst_i_2_n_0 ;
  wire \RD2_OBUF[2]_inst_i_3_n_0 ;
  wire \RD2_OBUF[2]_inst_i_4_n_0 ;
  wire \RD2_OBUF[2]_inst_i_5_n_0 ;
  wire \RD2_OBUF[2]_inst_i_6_n_0 ;
  wire \RD2_OBUF[2]_inst_i_7_n_0 ;
  wire \RD2_OBUF[2]_inst_i_8_n_0 ;
  wire \RD2_OBUF[2]_inst_i_9_n_0 ;
  wire \RD2_OBUF[30]_inst_i_10_n_0 ;
  wire \RD2_OBUF[30]_inst_i_11_n_0 ;
  wire \RD2_OBUF[30]_inst_i_12_n_0 ;
  wire \RD2_OBUF[30]_inst_i_13_n_0 ;
  wire \RD2_OBUF[30]_inst_i_2_n_0 ;
  wire \RD2_OBUF[30]_inst_i_3_n_0 ;
  wire \RD2_OBUF[30]_inst_i_4_n_0 ;
  wire \RD2_OBUF[30]_inst_i_5_n_0 ;
  wire \RD2_OBUF[30]_inst_i_6_n_0 ;
  wire \RD2_OBUF[30]_inst_i_7_n_0 ;
  wire \RD2_OBUF[30]_inst_i_8_n_0 ;
  wire \RD2_OBUF[30]_inst_i_9_n_0 ;
  wire \RD2_OBUF[31]_inst_i_10_n_0 ;
  wire \RD2_OBUF[31]_inst_i_11_n_0 ;
  wire \RD2_OBUF[31]_inst_i_12_n_0 ;
  wire \RD2_OBUF[31]_inst_i_13_n_0 ;
  wire \RD2_OBUF[31]_inst_i_2_n_0 ;
  wire \RD2_OBUF[31]_inst_i_3_n_0 ;
  wire \RD2_OBUF[31]_inst_i_4_n_0 ;
  wire \RD2_OBUF[31]_inst_i_5_n_0 ;
  wire \RD2_OBUF[31]_inst_i_6_n_0 ;
  wire \RD2_OBUF[31]_inst_i_7_n_0 ;
  wire \RD2_OBUF[31]_inst_i_8_n_0 ;
  wire \RD2_OBUF[31]_inst_i_9_n_0 ;
  wire \RD2_OBUF[3]_inst_i_10_n_0 ;
  wire \RD2_OBUF[3]_inst_i_11_n_0 ;
  wire \RD2_OBUF[3]_inst_i_12_n_0 ;
  wire \RD2_OBUF[3]_inst_i_13_n_0 ;
  wire \RD2_OBUF[3]_inst_i_2_n_0 ;
  wire \RD2_OBUF[3]_inst_i_3_n_0 ;
  wire \RD2_OBUF[3]_inst_i_4_n_0 ;
  wire \RD2_OBUF[3]_inst_i_5_n_0 ;
  wire \RD2_OBUF[3]_inst_i_6_n_0 ;
  wire \RD2_OBUF[3]_inst_i_7_n_0 ;
  wire \RD2_OBUF[3]_inst_i_8_n_0 ;
  wire \RD2_OBUF[3]_inst_i_9_n_0 ;
  wire \RD2_OBUF[4]_inst_i_10_n_0 ;
  wire \RD2_OBUF[4]_inst_i_11_n_0 ;
  wire \RD2_OBUF[4]_inst_i_12_n_0 ;
  wire \RD2_OBUF[4]_inst_i_13_n_0 ;
  wire \RD2_OBUF[4]_inst_i_2_n_0 ;
  wire \RD2_OBUF[4]_inst_i_3_n_0 ;
  wire \RD2_OBUF[4]_inst_i_4_n_0 ;
  wire \RD2_OBUF[4]_inst_i_5_n_0 ;
  wire \RD2_OBUF[4]_inst_i_6_n_0 ;
  wire \RD2_OBUF[4]_inst_i_7_n_0 ;
  wire \RD2_OBUF[4]_inst_i_8_n_0 ;
  wire \RD2_OBUF[4]_inst_i_9_n_0 ;
  wire \RD2_OBUF[5]_inst_i_10_n_0 ;
  wire \RD2_OBUF[5]_inst_i_11_n_0 ;
  wire \RD2_OBUF[5]_inst_i_12_n_0 ;
  wire \RD2_OBUF[5]_inst_i_13_n_0 ;
  wire \RD2_OBUF[5]_inst_i_2_n_0 ;
  wire \RD2_OBUF[5]_inst_i_3_n_0 ;
  wire \RD2_OBUF[5]_inst_i_4_n_0 ;
  wire \RD2_OBUF[5]_inst_i_5_n_0 ;
  wire \RD2_OBUF[5]_inst_i_6_n_0 ;
  wire \RD2_OBUF[5]_inst_i_7_n_0 ;
  wire \RD2_OBUF[5]_inst_i_8_n_0 ;
  wire \RD2_OBUF[5]_inst_i_9_n_0 ;
  wire \RD2_OBUF[6]_inst_i_10_n_0 ;
  wire \RD2_OBUF[6]_inst_i_11_n_0 ;
  wire \RD2_OBUF[6]_inst_i_12_n_0 ;
  wire \RD2_OBUF[6]_inst_i_13_n_0 ;
  wire \RD2_OBUF[6]_inst_i_2_n_0 ;
  wire \RD2_OBUF[6]_inst_i_3_n_0 ;
  wire \RD2_OBUF[6]_inst_i_4_n_0 ;
  wire \RD2_OBUF[6]_inst_i_5_n_0 ;
  wire \RD2_OBUF[6]_inst_i_6_n_0 ;
  wire \RD2_OBUF[6]_inst_i_7_n_0 ;
  wire \RD2_OBUF[6]_inst_i_8_n_0 ;
  wire \RD2_OBUF[6]_inst_i_9_n_0 ;
  wire \RD2_OBUF[7]_inst_i_10_n_0 ;
  wire \RD2_OBUF[7]_inst_i_11_n_0 ;
  wire \RD2_OBUF[7]_inst_i_12_n_0 ;
  wire \RD2_OBUF[7]_inst_i_13_n_0 ;
  wire \RD2_OBUF[7]_inst_i_2_n_0 ;
  wire \RD2_OBUF[7]_inst_i_3_n_0 ;
  wire \RD2_OBUF[7]_inst_i_4_n_0 ;
  wire \RD2_OBUF[7]_inst_i_5_n_0 ;
  wire \RD2_OBUF[7]_inst_i_6_n_0 ;
  wire \RD2_OBUF[7]_inst_i_7_n_0 ;
  wire \RD2_OBUF[7]_inst_i_8_n_0 ;
  wire \RD2_OBUF[7]_inst_i_9_n_0 ;
  wire \RD2_OBUF[8]_inst_i_10_n_0 ;
  wire \RD2_OBUF[8]_inst_i_11_n_0 ;
  wire \RD2_OBUF[8]_inst_i_12_n_0 ;
  wire \RD2_OBUF[8]_inst_i_13_n_0 ;
  wire \RD2_OBUF[8]_inst_i_2_n_0 ;
  wire \RD2_OBUF[8]_inst_i_3_n_0 ;
  wire \RD2_OBUF[8]_inst_i_4_n_0 ;
  wire \RD2_OBUF[8]_inst_i_5_n_0 ;
  wire \RD2_OBUF[8]_inst_i_6_n_0 ;
  wire \RD2_OBUF[8]_inst_i_7_n_0 ;
  wire \RD2_OBUF[8]_inst_i_8_n_0 ;
  wire \RD2_OBUF[8]_inst_i_9_n_0 ;
  wire \RD2_OBUF[9]_inst_i_10_n_0 ;
  wire \RD2_OBUF[9]_inst_i_11_n_0 ;
  wire \RD2_OBUF[9]_inst_i_12_n_0 ;
  wire \RD2_OBUF[9]_inst_i_13_n_0 ;
  wire \RD2_OBUF[9]_inst_i_2_n_0 ;
  wire \RD2_OBUF[9]_inst_i_3_n_0 ;
  wire \RD2_OBUF[9]_inst_i_4_n_0 ;
  wire \RD2_OBUF[9]_inst_i_5_n_0 ;
  wire \RD2_OBUF[9]_inst_i_6_n_0 ;
  wire \RD2_OBUF[9]_inst_i_7_n_0 ;
  wire \RD2_OBUF[9]_inst_i_8_n_0 ;
  wire \RD2_OBUF[9]_inst_i_9_n_0 ;
  wire [31:0]WD;
  wire [31:0]WD_IBUF;
  wire WE;
  wire WE_IBUF;
  wire clk;
  wire clk_IBUF;
  wire clk_IBUF_BUFG;
  wire r1;
  wire r10;
  wire \r10_reg_n_0_[0] ;
  wire \r10_reg_n_0_[10] ;
  wire \r10_reg_n_0_[11] ;
  wire \r10_reg_n_0_[12] ;
  wire \r10_reg_n_0_[13] ;
  wire \r10_reg_n_0_[14] ;
  wire \r10_reg_n_0_[15] ;
  wire \r10_reg_n_0_[16] ;
  wire \r10_reg_n_0_[17] ;
  wire \r10_reg_n_0_[18] ;
  wire \r10_reg_n_0_[19] ;
  wire \r10_reg_n_0_[1] ;
  wire \r10_reg_n_0_[20] ;
  wire \r10_reg_n_0_[21] ;
  wire \r10_reg_n_0_[22] ;
  wire \r10_reg_n_0_[23] ;
  wire \r10_reg_n_0_[24] ;
  wire \r10_reg_n_0_[25] ;
  wire \r10_reg_n_0_[26] ;
  wire \r10_reg_n_0_[27] ;
  wire \r10_reg_n_0_[28] ;
  wire \r10_reg_n_0_[29] ;
  wire \r10_reg_n_0_[2] ;
  wire \r10_reg_n_0_[30] ;
  wire \r10_reg_n_0_[31] ;
  wire \r10_reg_n_0_[3] ;
  wire \r10_reg_n_0_[4] ;
  wire \r10_reg_n_0_[5] ;
  wire \r10_reg_n_0_[6] ;
  wire \r10_reg_n_0_[7] ;
  wire \r10_reg_n_0_[8] ;
  wire \r10_reg_n_0_[9] ;
  wire r11;
  wire \r11_reg_n_0_[0] ;
  wire \r11_reg_n_0_[10] ;
  wire \r11_reg_n_0_[11] ;
  wire \r11_reg_n_0_[12] ;
  wire \r11_reg_n_0_[13] ;
  wire \r11_reg_n_0_[14] ;
  wire \r11_reg_n_0_[15] ;
  wire \r11_reg_n_0_[16] ;
  wire \r11_reg_n_0_[17] ;
  wire \r11_reg_n_0_[18] ;
  wire \r11_reg_n_0_[19] ;
  wire \r11_reg_n_0_[1] ;
  wire \r11_reg_n_0_[20] ;
  wire \r11_reg_n_0_[21] ;
  wire \r11_reg_n_0_[22] ;
  wire \r11_reg_n_0_[23] ;
  wire \r11_reg_n_0_[24] ;
  wire \r11_reg_n_0_[25] ;
  wire \r11_reg_n_0_[26] ;
  wire \r11_reg_n_0_[27] ;
  wire \r11_reg_n_0_[28] ;
  wire \r11_reg_n_0_[29] ;
  wire \r11_reg_n_0_[2] ;
  wire \r11_reg_n_0_[30] ;
  wire \r11_reg_n_0_[31] ;
  wire \r11_reg_n_0_[3] ;
  wire \r11_reg_n_0_[4] ;
  wire \r11_reg_n_0_[5] ;
  wire \r11_reg_n_0_[6] ;
  wire \r11_reg_n_0_[7] ;
  wire \r11_reg_n_0_[8] ;
  wire \r11_reg_n_0_[9] ;
  wire r12;
  wire \r12_reg_n_0_[0] ;
  wire \r12_reg_n_0_[10] ;
  wire \r12_reg_n_0_[11] ;
  wire \r12_reg_n_0_[12] ;
  wire \r12_reg_n_0_[13] ;
  wire \r12_reg_n_0_[14] ;
  wire \r12_reg_n_0_[15] ;
  wire \r12_reg_n_0_[16] ;
  wire \r12_reg_n_0_[17] ;
  wire \r12_reg_n_0_[18] ;
  wire \r12_reg_n_0_[19] ;
  wire \r12_reg_n_0_[1] ;
  wire \r12_reg_n_0_[20] ;
  wire \r12_reg_n_0_[21] ;
  wire \r12_reg_n_0_[22] ;
  wire \r12_reg_n_0_[23] ;
  wire \r12_reg_n_0_[24] ;
  wire \r12_reg_n_0_[25] ;
  wire \r12_reg_n_0_[26] ;
  wire \r12_reg_n_0_[27] ;
  wire \r12_reg_n_0_[28] ;
  wire \r12_reg_n_0_[29] ;
  wire \r12_reg_n_0_[2] ;
  wire \r12_reg_n_0_[30] ;
  wire \r12_reg_n_0_[31] ;
  wire \r12_reg_n_0_[3] ;
  wire \r12_reg_n_0_[4] ;
  wire \r12_reg_n_0_[5] ;
  wire \r12_reg_n_0_[6] ;
  wire \r12_reg_n_0_[7] ;
  wire \r12_reg_n_0_[8] ;
  wire \r12_reg_n_0_[9] ;
  wire r13;
  wire \r13_reg_n_0_[0] ;
  wire \r13_reg_n_0_[10] ;
  wire \r13_reg_n_0_[11] ;
  wire \r13_reg_n_0_[12] ;
  wire \r13_reg_n_0_[13] ;
  wire \r13_reg_n_0_[14] ;
  wire \r13_reg_n_0_[15] ;
  wire \r13_reg_n_0_[16] ;
  wire \r13_reg_n_0_[17] ;
  wire \r13_reg_n_0_[18] ;
  wire \r13_reg_n_0_[19] ;
  wire \r13_reg_n_0_[1] ;
  wire \r13_reg_n_0_[20] ;
  wire \r13_reg_n_0_[21] ;
  wire \r13_reg_n_0_[22] ;
  wire \r13_reg_n_0_[23] ;
  wire \r13_reg_n_0_[24] ;
  wire \r13_reg_n_0_[25] ;
  wire \r13_reg_n_0_[26] ;
  wire \r13_reg_n_0_[27] ;
  wire \r13_reg_n_0_[28] ;
  wire \r13_reg_n_0_[29] ;
  wire \r13_reg_n_0_[2] ;
  wire \r13_reg_n_0_[30] ;
  wire \r13_reg_n_0_[31] ;
  wire \r13_reg_n_0_[3] ;
  wire \r13_reg_n_0_[4] ;
  wire \r13_reg_n_0_[5] ;
  wire \r13_reg_n_0_[6] ;
  wire \r13_reg_n_0_[7] ;
  wire \r13_reg_n_0_[8] ;
  wire \r13_reg_n_0_[9] ;
  wire r14;
  wire \r14_reg_n_0_[0] ;
  wire \r14_reg_n_0_[10] ;
  wire \r14_reg_n_0_[11] ;
  wire \r14_reg_n_0_[12] ;
  wire \r14_reg_n_0_[13] ;
  wire \r14_reg_n_0_[14] ;
  wire \r14_reg_n_0_[15] ;
  wire \r14_reg_n_0_[16] ;
  wire \r14_reg_n_0_[17] ;
  wire \r14_reg_n_0_[18] ;
  wire \r14_reg_n_0_[19] ;
  wire \r14_reg_n_0_[1] ;
  wire \r14_reg_n_0_[20] ;
  wire \r14_reg_n_0_[21] ;
  wire \r14_reg_n_0_[22] ;
  wire \r14_reg_n_0_[23] ;
  wire \r14_reg_n_0_[24] ;
  wire \r14_reg_n_0_[25] ;
  wire \r14_reg_n_0_[26] ;
  wire \r14_reg_n_0_[27] ;
  wire \r14_reg_n_0_[28] ;
  wire \r14_reg_n_0_[29] ;
  wire \r14_reg_n_0_[2] ;
  wire \r14_reg_n_0_[30] ;
  wire \r14_reg_n_0_[31] ;
  wire \r14_reg_n_0_[3] ;
  wire \r14_reg_n_0_[4] ;
  wire \r14_reg_n_0_[5] ;
  wire \r14_reg_n_0_[6] ;
  wire \r14_reg_n_0_[7] ;
  wire \r14_reg_n_0_[8] ;
  wire \r14_reg_n_0_[9] ;
  wire r15;
  wire \r15_reg_n_0_[0] ;
  wire \r15_reg_n_0_[10] ;
  wire \r15_reg_n_0_[11] ;
  wire \r15_reg_n_0_[12] ;
  wire \r15_reg_n_0_[13] ;
  wire \r15_reg_n_0_[14] ;
  wire \r15_reg_n_0_[15] ;
  wire \r15_reg_n_0_[16] ;
  wire \r15_reg_n_0_[17] ;
  wire \r15_reg_n_0_[18] ;
  wire \r15_reg_n_0_[19] ;
  wire \r15_reg_n_0_[1] ;
  wire \r15_reg_n_0_[20] ;
  wire \r15_reg_n_0_[21] ;
  wire \r15_reg_n_0_[22] ;
  wire \r15_reg_n_0_[23] ;
  wire \r15_reg_n_0_[24] ;
  wire \r15_reg_n_0_[25] ;
  wire \r15_reg_n_0_[26] ;
  wire \r15_reg_n_0_[27] ;
  wire \r15_reg_n_0_[28] ;
  wire \r15_reg_n_0_[29] ;
  wire \r15_reg_n_0_[2] ;
  wire \r15_reg_n_0_[30] ;
  wire \r15_reg_n_0_[31] ;
  wire \r15_reg_n_0_[3] ;
  wire \r15_reg_n_0_[4] ;
  wire \r15_reg_n_0_[5] ;
  wire \r15_reg_n_0_[6] ;
  wire \r15_reg_n_0_[7] ;
  wire \r15_reg_n_0_[8] ;
  wire \r15_reg_n_0_[9] ;
  wire r16;
  wire \r16_reg_n_0_[0] ;
  wire \r16_reg_n_0_[10] ;
  wire \r16_reg_n_0_[11] ;
  wire \r16_reg_n_0_[12] ;
  wire \r16_reg_n_0_[13] ;
  wire \r16_reg_n_0_[14] ;
  wire \r16_reg_n_0_[15] ;
  wire \r16_reg_n_0_[16] ;
  wire \r16_reg_n_0_[17] ;
  wire \r16_reg_n_0_[18] ;
  wire \r16_reg_n_0_[19] ;
  wire \r16_reg_n_0_[1] ;
  wire \r16_reg_n_0_[20] ;
  wire \r16_reg_n_0_[21] ;
  wire \r16_reg_n_0_[22] ;
  wire \r16_reg_n_0_[23] ;
  wire \r16_reg_n_0_[24] ;
  wire \r16_reg_n_0_[25] ;
  wire \r16_reg_n_0_[26] ;
  wire \r16_reg_n_0_[27] ;
  wire \r16_reg_n_0_[28] ;
  wire \r16_reg_n_0_[29] ;
  wire \r16_reg_n_0_[2] ;
  wire \r16_reg_n_0_[30] ;
  wire \r16_reg_n_0_[31] ;
  wire \r16_reg_n_0_[3] ;
  wire \r16_reg_n_0_[4] ;
  wire \r16_reg_n_0_[5] ;
  wire \r16_reg_n_0_[6] ;
  wire \r16_reg_n_0_[7] ;
  wire \r16_reg_n_0_[8] ;
  wire \r16_reg_n_0_[9] ;
  wire r17;
  wire \r17_reg_n_0_[0] ;
  wire \r17_reg_n_0_[10] ;
  wire \r17_reg_n_0_[11] ;
  wire \r17_reg_n_0_[12] ;
  wire \r17_reg_n_0_[13] ;
  wire \r17_reg_n_0_[14] ;
  wire \r17_reg_n_0_[15] ;
  wire \r17_reg_n_0_[16] ;
  wire \r17_reg_n_0_[17] ;
  wire \r17_reg_n_0_[18] ;
  wire \r17_reg_n_0_[19] ;
  wire \r17_reg_n_0_[1] ;
  wire \r17_reg_n_0_[20] ;
  wire \r17_reg_n_0_[21] ;
  wire \r17_reg_n_0_[22] ;
  wire \r17_reg_n_0_[23] ;
  wire \r17_reg_n_0_[24] ;
  wire \r17_reg_n_0_[25] ;
  wire \r17_reg_n_0_[26] ;
  wire \r17_reg_n_0_[27] ;
  wire \r17_reg_n_0_[28] ;
  wire \r17_reg_n_0_[29] ;
  wire \r17_reg_n_0_[2] ;
  wire \r17_reg_n_0_[30] ;
  wire \r17_reg_n_0_[31] ;
  wire \r17_reg_n_0_[3] ;
  wire \r17_reg_n_0_[4] ;
  wire \r17_reg_n_0_[5] ;
  wire \r17_reg_n_0_[6] ;
  wire \r17_reg_n_0_[7] ;
  wire \r17_reg_n_0_[8] ;
  wire \r17_reg_n_0_[9] ;
  wire r18;
  wire \r18_reg_n_0_[0] ;
  wire \r18_reg_n_0_[10] ;
  wire \r18_reg_n_0_[11] ;
  wire \r18_reg_n_0_[12] ;
  wire \r18_reg_n_0_[13] ;
  wire \r18_reg_n_0_[14] ;
  wire \r18_reg_n_0_[15] ;
  wire \r18_reg_n_0_[16] ;
  wire \r18_reg_n_0_[17] ;
  wire \r18_reg_n_0_[18] ;
  wire \r18_reg_n_0_[19] ;
  wire \r18_reg_n_0_[1] ;
  wire \r18_reg_n_0_[20] ;
  wire \r18_reg_n_0_[21] ;
  wire \r18_reg_n_0_[22] ;
  wire \r18_reg_n_0_[23] ;
  wire \r18_reg_n_0_[24] ;
  wire \r18_reg_n_0_[25] ;
  wire \r18_reg_n_0_[26] ;
  wire \r18_reg_n_0_[27] ;
  wire \r18_reg_n_0_[28] ;
  wire \r18_reg_n_0_[29] ;
  wire \r18_reg_n_0_[2] ;
  wire \r18_reg_n_0_[30] ;
  wire \r18_reg_n_0_[31] ;
  wire \r18_reg_n_0_[3] ;
  wire \r18_reg_n_0_[4] ;
  wire \r18_reg_n_0_[5] ;
  wire \r18_reg_n_0_[6] ;
  wire \r18_reg_n_0_[7] ;
  wire \r18_reg_n_0_[8] ;
  wire \r18_reg_n_0_[9] ;
  wire r19;
  wire \r19_reg_n_0_[0] ;
  wire \r19_reg_n_0_[10] ;
  wire \r19_reg_n_0_[11] ;
  wire \r19_reg_n_0_[12] ;
  wire \r19_reg_n_0_[13] ;
  wire \r19_reg_n_0_[14] ;
  wire \r19_reg_n_0_[15] ;
  wire \r19_reg_n_0_[16] ;
  wire \r19_reg_n_0_[17] ;
  wire \r19_reg_n_0_[18] ;
  wire \r19_reg_n_0_[19] ;
  wire \r19_reg_n_0_[1] ;
  wire \r19_reg_n_0_[20] ;
  wire \r19_reg_n_0_[21] ;
  wire \r19_reg_n_0_[22] ;
  wire \r19_reg_n_0_[23] ;
  wire \r19_reg_n_0_[24] ;
  wire \r19_reg_n_0_[25] ;
  wire \r19_reg_n_0_[26] ;
  wire \r19_reg_n_0_[27] ;
  wire \r19_reg_n_0_[28] ;
  wire \r19_reg_n_0_[29] ;
  wire \r19_reg_n_0_[2] ;
  wire \r19_reg_n_0_[30] ;
  wire \r19_reg_n_0_[31] ;
  wire \r19_reg_n_0_[3] ;
  wire \r19_reg_n_0_[4] ;
  wire \r19_reg_n_0_[5] ;
  wire \r19_reg_n_0_[6] ;
  wire \r19_reg_n_0_[7] ;
  wire \r19_reg_n_0_[8] ;
  wire \r19_reg_n_0_[9] ;
  wire \r1_reg_n_0_[0] ;
  wire \r1_reg_n_0_[10] ;
  wire \r1_reg_n_0_[11] ;
  wire \r1_reg_n_0_[12] ;
  wire \r1_reg_n_0_[13] ;
  wire \r1_reg_n_0_[14] ;
  wire \r1_reg_n_0_[15] ;
  wire \r1_reg_n_0_[16] ;
  wire \r1_reg_n_0_[17] ;
  wire \r1_reg_n_0_[18] ;
  wire \r1_reg_n_0_[19] ;
  wire \r1_reg_n_0_[1] ;
  wire \r1_reg_n_0_[20] ;
  wire \r1_reg_n_0_[21] ;
  wire \r1_reg_n_0_[22] ;
  wire \r1_reg_n_0_[23] ;
  wire \r1_reg_n_0_[24] ;
  wire \r1_reg_n_0_[25] ;
  wire \r1_reg_n_0_[26] ;
  wire \r1_reg_n_0_[27] ;
  wire \r1_reg_n_0_[28] ;
  wire \r1_reg_n_0_[29] ;
  wire \r1_reg_n_0_[2] ;
  wire \r1_reg_n_0_[30] ;
  wire \r1_reg_n_0_[31] ;
  wire \r1_reg_n_0_[3] ;
  wire \r1_reg_n_0_[4] ;
  wire \r1_reg_n_0_[5] ;
  wire \r1_reg_n_0_[6] ;
  wire \r1_reg_n_0_[7] ;
  wire \r1_reg_n_0_[8] ;
  wire \r1_reg_n_0_[9] ;
  wire r2;
  wire r20;
  wire \r20_reg_n_0_[0] ;
  wire \r20_reg_n_0_[10] ;
  wire \r20_reg_n_0_[11] ;
  wire \r20_reg_n_0_[12] ;
  wire \r20_reg_n_0_[13] ;
  wire \r20_reg_n_0_[14] ;
  wire \r20_reg_n_0_[15] ;
  wire \r20_reg_n_0_[16] ;
  wire \r20_reg_n_0_[17] ;
  wire \r20_reg_n_0_[18] ;
  wire \r20_reg_n_0_[19] ;
  wire \r20_reg_n_0_[1] ;
  wire \r20_reg_n_0_[20] ;
  wire \r20_reg_n_0_[21] ;
  wire \r20_reg_n_0_[22] ;
  wire \r20_reg_n_0_[23] ;
  wire \r20_reg_n_0_[24] ;
  wire \r20_reg_n_0_[25] ;
  wire \r20_reg_n_0_[26] ;
  wire \r20_reg_n_0_[27] ;
  wire \r20_reg_n_0_[28] ;
  wire \r20_reg_n_0_[29] ;
  wire \r20_reg_n_0_[2] ;
  wire \r20_reg_n_0_[30] ;
  wire \r20_reg_n_0_[31] ;
  wire \r20_reg_n_0_[3] ;
  wire \r20_reg_n_0_[4] ;
  wire \r20_reg_n_0_[5] ;
  wire \r20_reg_n_0_[6] ;
  wire \r20_reg_n_0_[7] ;
  wire \r20_reg_n_0_[8] ;
  wire \r20_reg_n_0_[9] ;
  wire r21;
  wire \r21_reg_n_0_[0] ;
  wire \r21_reg_n_0_[10] ;
  wire \r21_reg_n_0_[11] ;
  wire \r21_reg_n_0_[12] ;
  wire \r21_reg_n_0_[13] ;
  wire \r21_reg_n_0_[14] ;
  wire \r21_reg_n_0_[15] ;
  wire \r21_reg_n_0_[16] ;
  wire \r21_reg_n_0_[17] ;
  wire \r21_reg_n_0_[18] ;
  wire \r21_reg_n_0_[19] ;
  wire \r21_reg_n_0_[1] ;
  wire \r21_reg_n_0_[20] ;
  wire \r21_reg_n_0_[21] ;
  wire \r21_reg_n_0_[22] ;
  wire \r21_reg_n_0_[23] ;
  wire \r21_reg_n_0_[24] ;
  wire \r21_reg_n_0_[25] ;
  wire \r21_reg_n_0_[26] ;
  wire \r21_reg_n_0_[27] ;
  wire \r21_reg_n_0_[28] ;
  wire \r21_reg_n_0_[29] ;
  wire \r21_reg_n_0_[2] ;
  wire \r21_reg_n_0_[30] ;
  wire \r21_reg_n_0_[31] ;
  wire \r21_reg_n_0_[3] ;
  wire \r21_reg_n_0_[4] ;
  wire \r21_reg_n_0_[5] ;
  wire \r21_reg_n_0_[6] ;
  wire \r21_reg_n_0_[7] ;
  wire \r21_reg_n_0_[8] ;
  wire \r21_reg_n_0_[9] ;
  wire r22;
  wire \r22_reg_n_0_[0] ;
  wire \r22_reg_n_0_[10] ;
  wire \r22_reg_n_0_[11] ;
  wire \r22_reg_n_0_[12] ;
  wire \r22_reg_n_0_[13] ;
  wire \r22_reg_n_0_[14] ;
  wire \r22_reg_n_0_[15] ;
  wire \r22_reg_n_0_[16] ;
  wire \r22_reg_n_0_[17] ;
  wire \r22_reg_n_0_[18] ;
  wire \r22_reg_n_0_[19] ;
  wire \r22_reg_n_0_[1] ;
  wire \r22_reg_n_0_[20] ;
  wire \r22_reg_n_0_[21] ;
  wire \r22_reg_n_0_[22] ;
  wire \r22_reg_n_0_[23] ;
  wire \r22_reg_n_0_[24] ;
  wire \r22_reg_n_0_[25] ;
  wire \r22_reg_n_0_[26] ;
  wire \r22_reg_n_0_[27] ;
  wire \r22_reg_n_0_[28] ;
  wire \r22_reg_n_0_[29] ;
  wire \r22_reg_n_0_[2] ;
  wire \r22_reg_n_0_[30] ;
  wire \r22_reg_n_0_[31] ;
  wire \r22_reg_n_0_[3] ;
  wire \r22_reg_n_0_[4] ;
  wire \r22_reg_n_0_[5] ;
  wire \r22_reg_n_0_[6] ;
  wire \r22_reg_n_0_[7] ;
  wire \r22_reg_n_0_[8] ;
  wire \r22_reg_n_0_[9] ;
  wire r23;
  wire \r23_reg_n_0_[0] ;
  wire \r23_reg_n_0_[10] ;
  wire \r23_reg_n_0_[11] ;
  wire \r23_reg_n_0_[12] ;
  wire \r23_reg_n_0_[13] ;
  wire \r23_reg_n_0_[14] ;
  wire \r23_reg_n_0_[15] ;
  wire \r23_reg_n_0_[16] ;
  wire \r23_reg_n_0_[17] ;
  wire \r23_reg_n_0_[18] ;
  wire \r23_reg_n_0_[19] ;
  wire \r23_reg_n_0_[1] ;
  wire \r23_reg_n_0_[20] ;
  wire \r23_reg_n_0_[21] ;
  wire \r23_reg_n_0_[22] ;
  wire \r23_reg_n_0_[23] ;
  wire \r23_reg_n_0_[24] ;
  wire \r23_reg_n_0_[25] ;
  wire \r23_reg_n_0_[26] ;
  wire \r23_reg_n_0_[27] ;
  wire \r23_reg_n_0_[28] ;
  wire \r23_reg_n_0_[29] ;
  wire \r23_reg_n_0_[2] ;
  wire \r23_reg_n_0_[30] ;
  wire \r23_reg_n_0_[31] ;
  wire \r23_reg_n_0_[3] ;
  wire \r23_reg_n_0_[4] ;
  wire \r23_reg_n_0_[5] ;
  wire \r23_reg_n_0_[6] ;
  wire \r23_reg_n_0_[7] ;
  wire \r23_reg_n_0_[8] ;
  wire \r23_reg_n_0_[9] ;
  wire r24;
  wire \r24_reg_n_0_[0] ;
  wire \r24_reg_n_0_[10] ;
  wire \r24_reg_n_0_[11] ;
  wire \r24_reg_n_0_[12] ;
  wire \r24_reg_n_0_[13] ;
  wire \r24_reg_n_0_[14] ;
  wire \r24_reg_n_0_[15] ;
  wire \r24_reg_n_0_[16] ;
  wire \r24_reg_n_0_[17] ;
  wire \r24_reg_n_0_[18] ;
  wire \r24_reg_n_0_[19] ;
  wire \r24_reg_n_0_[1] ;
  wire \r24_reg_n_0_[20] ;
  wire \r24_reg_n_0_[21] ;
  wire \r24_reg_n_0_[22] ;
  wire \r24_reg_n_0_[23] ;
  wire \r24_reg_n_0_[24] ;
  wire \r24_reg_n_0_[25] ;
  wire \r24_reg_n_0_[26] ;
  wire \r24_reg_n_0_[27] ;
  wire \r24_reg_n_0_[28] ;
  wire \r24_reg_n_0_[29] ;
  wire \r24_reg_n_0_[2] ;
  wire \r24_reg_n_0_[30] ;
  wire \r24_reg_n_0_[31] ;
  wire \r24_reg_n_0_[3] ;
  wire \r24_reg_n_0_[4] ;
  wire \r24_reg_n_0_[5] ;
  wire \r24_reg_n_0_[6] ;
  wire \r24_reg_n_0_[7] ;
  wire \r24_reg_n_0_[8] ;
  wire \r24_reg_n_0_[9] ;
  wire r25;
  wire \r25_reg_n_0_[0] ;
  wire \r25_reg_n_0_[10] ;
  wire \r25_reg_n_0_[11] ;
  wire \r25_reg_n_0_[12] ;
  wire \r25_reg_n_0_[13] ;
  wire \r25_reg_n_0_[14] ;
  wire \r25_reg_n_0_[15] ;
  wire \r25_reg_n_0_[16] ;
  wire \r25_reg_n_0_[17] ;
  wire \r25_reg_n_0_[18] ;
  wire \r25_reg_n_0_[19] ;
  wire \r25_reg_n_0_[1] ;
  wire \r25_reg_n_0_[20] ;
  wire \r25_reg_n_0_[21] ;
  wire \r25_reg_n_0_[22] ;
  wire \r25_reg_n_0_[23] ;
  wire \r25_reg_n_0_[24] ;
  wire \r25_reg_n_0_[25] ;
  wire \r25_reg_n_0_[26] ;
  wire \r25_reg_n_0_[27] ;
  wire \r25_reg_n_0_[28] ;
  wire \r25_reg_n_0_[29] ;
  wire \r25_reg_n_0_[2] ;
  wire \r25_reg_n_0_[30] ;
  wire \r25_reg_n_0_[31] ;
  wire \r25_reg_n_0_[3] ;
  wire \r25_reg_n_0_[4] ;
  wire \r25_reg_n_0_[5] ;
  wire \r25_reg_n_0_[6] ;
  wire \r25_reg_n_0_[7] ;
  wire \r25_reg_n_0_[8] ;
  wire \r25_reg_n_0_[9] ;
  wire r26;
  wire \r26_reg_n_0_[0] ;
  wire \r26_reg_n_0_[10] ;
  wire \r26_reg_n_0_[11] ;
  wire \r26_reg_n_0_[12] ;
  wire \r26_reg_n_0_[13] ;
  wire \r26_reg_n_0_[14] ;
  wire \r26_reg_n_0_[15] ;
  wire \r26_reg_n_0_[16] ;
  wire \r26_reg_n_0_[17] ;
  wire \r26_reg_n_0_[18] ;
  wire \r26_reg_n_0_[19] ;
  wire \r26_reg_n_0_[1] ;
  wire \r26_reg_n_0_[20] ;
  wire \r26_reg_n_0_[21] ;
  wire \r26_reg_n_0_[22] ;
  wire \r26_reg_n_0_[23] ;
  wire \r26_reg_n_0_[24] ;
  wire \r26_reg_n_0_[25] ;
  wire \r26_reg_n_0_[26] ;
  wire \r26_reg_n_0_[27] ;
  wire \r26_reg_n_0_[28] ;
  wire \r26_reg_n_0_[29] ;
  wire \r26_reg_n_0_[2] ;
  wire \r26_reg_n_0_[30] ;
  wire \r26_reg_n_0_[31] ;
  wire \r26_reg_n_0_[3] ;
  wire \r26_reg_n_0_[4] ;
  wire \r26_reg_n_0_[5] ;
  wire \r26_reg_n_0_[6] ;
  wire \r26_reg_n_0_[7] ;
  wire \r26_reg_n_0_[8] ;
  wire \r26_reg_n_0_[9] ;
  wire r27;
  wire \r27_reg_n_0_[0] ;
  wire \r27_reg_n_0_[10] ;
  wire \r27_reg_n_0_[11] ;
  wire \r27_reg_n_0_[12] ;
  wire \r27_reg_n_0_[13] ;
  wire \r27_reg_n_0_[14] ;
  wire \r27_reg_n_0_[15] ;
  wire \r27_reg_n_0_[16] ;
  wire \r27_reg_n_0_[17] ;
  wire \r27_reg_n_0_[18] ;
  wire \r27_reg_n_0_[19] ;
  wire \r27_reg_n_0_[1] ;
  wire \r27_reg_n_0_[20] ;
  wire \r27_reg_n_0_[21] ;
  wire \r27_reg_n_0_[22] ;
  wire \r27_reg_n_0_[23] ;
  wire \r27_reg_n_0_[24] ;
  wire \r27_reg_n_0_[25] ;
  wire \r27_reg_n_0_[26] ;
  wire \r27_reg_n_0_[27] ;
  wire \r27_reg_n_0_[28] ;
  wire \r27_reg_n_0_[29] ;
  wire \r27_reg_n_0_[2] ;
  wire \r27_reg_n_0_[30] ;
  wire \r27_reg_n_0_[31] ;
  wire \r27_reg_n_0_[3] ;
  wire \r27_reg_n_0_[4] ;
  wire \r27_reg_n_0_[5] ;
  wire \r27_reg_n_0_[6] ;
  wire \r27_reg_n_0_[7] ;
  wire \r27_reg_n_0_[8] ;
  wire \r27_reg_n_0_[9] ;
  wire r28;
  wire \r28_reg_n_0_[0] ;
  wire \r28_reg_n_0_[10] ;
  wire \r28_reg_n_0_[11] ;
  wire \r28_reg_n_0_[12] ;
  wire \r28_reg_n_0_[13] ;
  wire \r28_reg_n_0_[14] ;
  wire \r28_reg_n_0_[15] ;
  wire \r28_reg_n_0_[16] ;
  wire \r28_reg_n_0_[17] ;
  wire \r28_reg_n_0_[18] ;
  wire \r28_reg_n_0_[19] ;
  wire \r28_reg_n_0_[1] ;
  wire \r28_reg_n_0_[20] ;
  wire \r28_reg_n_0_[21] ;
  wire \r28_reg_n_0_[22] ;
  wire \r28_reg_n_0_[23] ;
  wire \r28_reg_n_0_[24] ;
  wire \r28_reg_n_0_[25] ;
  wire \r28_reg_n_0_[26] ;
  wire \r28_reg_n_0_[27] ;
  wire \r28_reg_n_0_[28] ;
  wire \r28_reg_n_0_[29] ;
  wire \r28_reg_n_0_[2] ;
  wire \r28_reg_n_0_[30] ;
  wire \r28_reg_n_0_[31] ;
  wire \r28_reg_n_0_[3] ;
  wire \r28_reg_n_0_[4] ;
  wire \r28_reg_n_0_[5] ;
  wire \r28_reg_n_0_[6] ;
  wire \r28_reg_n_0_[7] ;
  wire \r28_reg_n_0_[8] ;
  wire \r28_reg_n_0_[9] ;
  wire r29;
  wire \r29_reg_n_0_[0] ;
  wire \r29_reg_n_0_[10] ;
  wire \r29_reg_n_0_[11] ;
  wire \r29_reg_n_0_[12] ;
  wire \r29_reg_n_0_[13] ;
  wire \r29_reg_n_0_[14] ;
  wire \r29_reg_n_0_[15] ;
  wire \r29_reg_n_0_[16] ;
  wire \r29_reg_n_0_[17] ;
  wire \r29_reg_n_0_[18] ;
  wire \r29_reg_n_0_[19] ;
  wire \r29_reg_n_0_[1] ;
  wire \r29_reg_n_0_[20] ;
  wire \r29_reg_n_0_[21] ;
  wire \r29_reg_n_0_[22] ;
  wire \r29_reg_n_0_[23] ;
  wire \r29_reg_n_0_[24] ;
  wire \r29_reg_n_0_[25] ;
  wire \r29_reg_n_0_[26] ;
  wire \r29_reg_n_0_[27] ;
  wire \r29_reg_n_0_[28] ;
  wire \r29_reg_n_0_[29] ;
  wire \r29_reg_n_0_[2] ;
  wire \r29_reg_n_0_[30] ;
  wire \r29_reg_n_0_[31] ;
  wire \r29_reg_n_0_[3] ;
  wire \r29_reg_n_0_[4] ;
  wire \r29_reg_n_0_[5] ;
  wire \r29_reg_n_0_[6] ;
  wire \r29_reg_n_0_[7] ;
  wire \r29_reg_n_0_[8] ;
  wire \r29_reg_n_0_[9] ;
  wire \r2_reg_n_0_[0] ;
  wire \r2_reg_n_0_[10] ;
  wire \r2_reg_n_0_[11] ;
  wire \r2_reg_n_0_[12] ;
  wire \r2_reg_n_0_[13] ;
  wire \r2_reg_n_0_[14] ;
  wire \r2_reg_n_0_[15] ;
  wire \r2_reg_n_0_[16] ;
  wire \r2_reg_n_0_[17] ;
  wire \r2_reg_n_0_[18] ;
  wire \r2_reg_n_0_[19] ;
  wire \r2_reg_n_0_[1] ;
  wire \r2_reg_n_0_[20] ;
  wire \r2_reg_n_0_[21] ;
  wire \r2_reg_n_0_[22] ;
  wire \r2_reg_n_0_[23] ;
  wire \r2_reg_n_0_[24] ;
  wire \r2_reg_n_0_[25] ;
  wire \r2_reg_n_0_[26] ;
  wire \r2_reg_n_0_[27] ;
  wire \r2_reg_n_0_[28] ;
  wire \r2_reg_n_0_[29] ;
  wire \r2_reg_n_0_[2] ;
  wire \r2_reg_n_0_[30] ;
  wire \r2_reg_n_0_[31] ;
  wire \r2_reg_n_0_[3] ;
  wire \r2_reg_n_0_[4] ;
  wire \r2_reg_n_0_[5] ;
  wire \r2_reg_n_0_[6] ;
  wire \r2_reg_n_0_[7] ;
  wire \r2_reg_n_0_[8] ;
  wire \r2_reg_n_0_[9] ;
  wire r3;
  wire r30;
  wire \r30_reg_n_0_[0] ;
  wire \r30_reg_n_0_[10] ;
  wire \r30_reg_n_0_[11] ;
  wire \r30_reg_n_0_[12] ;
  wire \r30_reg_n_0_[13] ;
  wire \r30_reg_n_0_[14] ;
  wire \r30_reg_n_0_[15] ;
  wire \r30_reg_n_0_[16] ;
  wire \r30_reg_n_0_[17] ;
  wire \r30_reg_n_0_[18] ;
  wire \r30_reg_n_0_[19] ;
  wire \r30_reg_n_0_[1] ;
  wire \r30_reg_n_0_[20] ;
  wire \r30_reg_n_0_[21] ;
  wire \r30_reg_n_0_[22] ;
  wire \r30_reg_n_0_[23] ;
  wire \r30_reg_n_0_[24] ;
  wire \r30_reg_n_0_[25] ;
  wire \r30_reg_n_0_[26] ;
  wire \r30_reg_n_0_[27] ;
  wire \r30_reg_n_0_[28] ;
  wire \r30_reg_n_0_[29] ;
  wire \r30_reg_n_0_[2] ;
  wire \r30_reg_n_0_[30] ;
  wire \r30_reg_n_0_[31] ;
  wire \r30_reg_n_0_[3] ;
  wire \r30_reg_n_0_[4] ;
  wire \r30_reg_n_0_[5] ;
  wire \r30_reg_n_0_[6] ;
  wire \r30_reg_n_0_[7] ;
  wire \r30_reg_n_0_[8] ;
  wire \r30_reg_n_0_[9] ;
  wire r31;
  wire \r31_reg_n_0_[0] ;
  wire \r31_reg_n_0_[10] ;
  wire \r31_reg_n_0_[11] ;
  wire \r31_reg_n_0_[12] ;
  wire \r31_reg_n_0_[13] ;
  wire \r31_reg_n_0_[14] ;
  wire \r31_reg_n_0_[15] ;
  wire \r31_reg_n_0_[16] ;
  wire \r31_reg_n_0_[17] ;
  wire \r31_reg_n_0_[18] ;
  wire \r31_reg_n_0_[19] ;
  wire \r31_reg_n_0_[1] ;
  wire \r31_reg_n_0_[20] ;
  wire \r31_reg_n_0_[21] ;
  wire \r31_reg_n_0_[22] ;
  wire \r31_reg_n_0_[23] ;
  wire \r31_reg_n_0_[24] ;
  wire \r31_reg_n_0_[25] ;
  wire \r31_reg_n_0_[26] ;
  wire \r31_reg_n_0_[27] ;
  wire \r31_reg_n_0_[28] ;
  wire \r31_reg_n_0_[29] ;
  wire \r31_reg_n_0_[2] ;
  wire \r31_reg_n_0_[30] ;
  wire \r31_reg_n_0_[31] ;
  wire \r31_reg_n_0_[3] ;
  wire \r31_reg_n_0_[4] ;
  wire \r31_reg_n_0_[5] ;
  wire \r31_reg_n_0_[6] ;
  wire \r31_reg_n_0_[7] ;
  wire \r31_reg_n_0_[8] ;
  wire \r31_reg_n_0_[9] ;
  wire \r3_reg_n_0_[0] ;
  wire \r3_reg_n_0_[10] ;
  wire \r3_reg_n_0_[11] ;
  wire \r3_reg_n_0_[12] ;
  wire \r3_reg_n_0_[13] ;
  wire \r3_reg_n_0_[14] ;
  wire \r3_reg_n_0_[15] ;
  wire \r3_reg_n_0_[16] ;
  wire \r3_reg_n_0_[17] ;
  wire \r3_reg_n_0_[18] ;
  wire \r3_reg_n_0_[19] ;
  wire \r3_reg_n_0_[1] ;
  wire \r3_reg_n_0_[20] ;
  wire \r3_reg_n_0_[21] ;
  wire \r3_reg_n_0_[22] ;
  wire \r3_reg_n_0_[23] ;
  wire \r3_reg_n_0_[24] ;
  wire \r3_reg_n_0_[25] ;
  wire \r3_reg_n_0_[26] ;
  wire \r3_reg_n_0_[27] ;
  wire \r3_reg_n_0_[28] ;
  wire \r3_reg_n_0_[29] ;
  wire \r3_reg_n_0_[2] ;
  wire \r3_reg_n_0_[30] ;
  wire \r3_reg_n_0_[31] ;
  wire \r3_reg_n_0_[3] ;
  wire \r3_reg_n_0_[4] ;
  wire \r3_reg_n_0_[5] ;
  wire \r3_reg_n_0_[6] ;
  wire \r3_reg_n_0_[7] ;
  wire \r3_reg_n_0_[8] ;
  wire \r3_reg_n_0_[9] ;
  wire r4;
  wire \r4_reg_n_0_[0] ;
  wire \r4_reg_n_0_[10] ;
  wire \r4_reg_n_0_[11] ;
  wire \r4_reg_n_0_[12] ;
  wire \r4_reg_n_0_[13] ;
  wire \r4_reg_n_0_[14] ;
  wire \r4_reg_n_0_[15] ;
  wire \r4_reg_n_0_[16] ;
  wire \r4_reg_n_0_[17] ;
  wire \r4_reg_n_0_[18] ;
  wire \r4_reg_n_0_[19] ;
  wire \r4_reg_n_0_[1] ;
  wire \r4_reg_n_0_[20] ;
  wire \r4_reg_n_0_[21] ;
  wire \r4_reg_n_0_[22] ;
  wire \r4_reg_n_0_[23] ;
  wire \r4_reg_n_0_[24] ;
  wire \r4_reg_n_0_[25] ;
  wire \r4_reg_n_0_[26] ;
  wire \r4_reg_n_0_[27] ;
  wire \r4_reg_n_0_[28] ;
  wire \r4_reg_n_0_[29] ;
  wire \r4_reg_n_0_[2] ;
  wire \r4_reg_n_0_[30] ;
  wire \r4_reg_n_0_[31] ;
  wire \r4_reg_n_0_[3] ;
  wire \r4_reg_n_0_[4] ;
  wire \r4_reg_n_0_[5] ;
  wire \r4_reg_n_0_[6] ;
  wire \r4_reg_n_0_[7] ;
  wire \r4_reg_n_0_[8] ;
  wire \r4_reg_n_0_[9] ;
  wire r5;
  wire \r5_reg_n_0_[0] ;
  wire \r5_reg_n_0_[10] ;
  wire \r5_reg_n_0_[11] ;
  wire \r5_reg_n_0_[12] ;
  wire \r5_reg_n_0_[13] ;
  wire \r5_reg_n_0_[14] ;
  wire \r5_reg_n_0_[15] ;
  wire \r5_reg_n_0_[16] ;
  wire \r5_reg_n_0_[17] ;
  wire \r5_reg_n_0_[18] ;
  wire \r5_reg_n_0_[19] ;
  wire \r5_reg_n_0_[1] ;
  wire \r5_reg_n_0_[20] ;
  wire \r5_reg_n_0_[21] ;
  wire \r5_reg_n_0_[22] ;
  wire \r5_reg_n_0_[23] ;
  wire \r5_reg_n_0_[24] ;
  wire \r5_reg_n_0_[25] ;
  wire \r5_reg_n_0_[26] ;
  wire \r5_reg_n_0_[27] ;
  wire \r5_reg_n_0_[28] ;
  wire \r5_reg_n_0_[29] ;
  wire \r5_reg_n_0_[2] ;
  wire \r5_reg_n_0_[30] ;
  wire \r5_reg_n_0_[31] ;
  wire \r5_reg_n_0_[3] ;
  wire \r5_reg_n_0_[4] ;
  wire \r5_reg_n_0_[5] ;
  wire \r5_reg_n_0_[6] ;
  wire \r5_reg_n_0_[7] ;
  wire \r5_reg_n_0_[8] ;
  wire \r5_reg_n_0_[9] ;
  wire r6;
  wire \r6_reg_n_0_[0] ;
  wire \r6_reg_n_0_[10] ;
  wire \r6_reg_n_0_[11] ;
  wire \r6_reg_n_0_[12] ;
  wire \r6_reg_n_0_[13] ;
  wire \r6_reg_n_0_[14] ;
  wire \r6_reg_n_0_[15] ;
  wire \r6_reg_n_0_[16] ;
  wire \r6_reg_n_0_[17] ;
  wire \r6_reg_n_0_[18] ;
  wire \r6_reg_n_0_[19] ;
  wire \r6_reg_n_0_[1] ;
  wire \r6_reg_n_0_[20] ;
  wire \r6_reg_n_0_[21] ;
  wire \r6_reg_n_0_[22] ;
  wire \r6_reg_n_0_[23] ;
  wire \r6_reg_n_0_[24] ;
  wire \r6_reg_n_0_[25] ;
  wire \r6_reg_n_0_[26] ;
  wire \r6_reg_n_0_[27] ;
  wire \r6_reg_n_0_[28] ;
  wire \r6_reg_n_0_[29] ;
  wire \r6_reg_n_0_[2] ;
  wire \r6_reg_n_0_[30] ;
  wire \r6_reg_n_0_[31] ;
  wire \r6_reg_n_0_[3] ;
  wire \r6_reg_n_0_[4] ;
  wire \r6_reg_n_0_[5] ;
  wire \r6_reg_n_0_[6] ;
  wire \r6_reg_n_0_[7] ;
  wire \r6_reg_n_0_[8] ;
  wire \r6_reg_n_0_[9] ;
  wire r7;
  wire \r7_reg_n_0_[0] ;
  wire \r7_reg_n_0_[10] ;
  wire \r7_reg_n_0_[11] ;
  wire \r7_reg_n_0_[12] ;
  wire \r7_reg_n_0_[13] ;
  wire \r7_reg_n_0_[14] ;
  wire \r7_reg_n_0_[15] ;
  wire \r7_reg_n_0_[16] ;
  wire \r7_reg_n_0_[17] ;
  wire \r7_reg_n_0_[18] ;
  wire \r7_reg_n_0_[19] ;
  wire \r7_reg_n_0_[1] ;
  wire \r7_reg_n_0_[20] ;
  wire \r7_reg_n_0_[21] ;
  wire \r7_reg_n_0_[22] ;
  wire \r7_reg_n_0_[23] ;
  wire \r7_reg_n_0_[24] ;
  wire \r7_reg_n_0_[25] ;
  wire \r7_reg_n_0_[26] ;
  wire \r7_reg_n_0_[27] ;
  wire \r7_reg_n_0_[28] ;
  wire \r7_reg_n_0_[29] ;
  wire \r7_reg_n_0_[2] ;
  wire \r7_reg_n_0_[30] ;
  wire \r7_reg_n_0_[31] ;
  wire \r7_reg_n_0_[3] ;
  wire \r7_reg_n_0_[4] ;
  wire \r7_reg_n_0_[5] ;
  wire \r7_reg_n_0_[6] ;
  wire \r7_reg_n_0_[7] ;
  wire \r7_reg_n_0_[8] ;
  wire \r7_reg_n_0_[9] ;
  wire r8;
  wire \r8_reg_n_0_[0] ;
  wire \r8_reg_n_0_[10] ;
  wire \r8_reg_n_0_[11] ;
  wire \r8_reg_n_0_[12] ;
  wire \r8_reg_n_0_[13] ;
  wire \r8_reg_n_0_[14] ;
  wire \r8_reg_n_0_[15] ;
  wire \r8_reg_n_0_[16] ;
  wire \r8_reg_n_0_[17] ;
  wire \r8_reg_n_0_[18] ;
  wire \r8_reg_n_0_[19] ;
  wire \r8_reg_n_0_[1] ;
  wire \r8_reg_n_0_[20] ;
  wire \r8_reg_n_0_[21] ;
  wire \r8_reg_n_0_[22] ;
  wire \r8_reg_n_0_[23] ;
  wire \r8_reg_n_0_[24] ;
  wire \r8_reg_n_0_[25] ;
  wire \r8_reg_n_0_[26] ;
  wire \r8_reg_n_0_[27] ;
  wire \r8_reg_n_0_[28] ;
  wire \r8_reg_n_0_[29] ;
  wire \r8_reg_n_0_[2] ;
  wire \r8_reg_n_0_[30] ;
  wire \r8_reg_n_0_[31] ;
  wire \r8_reg_n_0_[3] ;
  wire \r8_reg_n_0_[4] ;
  wire \r8_reg_n_0_[5] ;
  wire \r8_reg_n_0_[6] ;
  wire \r8_reg_n_0_[7] ;
  wire \r8_reg_n_0_[8] ;
  wire \r8_reg_n_0_[9] ;
  wire r9;
  wire \r9_reg_n_0_[0] ;
  wire \r9_reg_n_0_[10] ;
  wire \r9_reg_n_0_[11] ;
  wire \r9_reg_n_0_[12] ;
  wire \r9_reg_n_0_[13] ;
  wire \r9_reg_n_0_[14] ;
  wire \r9_reg_n_0_[15] ;
  wire \r9_reg_n_0_[16] ;
  wire \r9_reg_n_0_[17] ;
  wire \r9_reg_n_0_[18] ;
  wire \r9_reg_n_0_[19] ;
  wire \r9_reg_n_0_[1] ;
  wire \r9_reg_n_0_[20] ;
  wire \r9_reg_n_0_[21] ;
  wire \r9_reg_n_0_[22] ;
  wire \r9_reg_n_0_[23] ;
  wire \r9_reg_n_0_[24] ;
  wire \r9_reg_n_0_[25] ;
  wire \r9_reg_n_0_[26] ;
  wire \r9_reg_n_0_[27] ;
  wire \r9_reg_n_0_[28] ;
  wire \r9_reg_n_0_[29] ;
  wire \r9_reg_n_0_[2] ;
  wire \r9_reg_n_0_[30] ;
  wire \r9_reg_n_0_[31] ;
  wire \r9_reg_n_0_[3] ;
  wire \r9_reg_n_0_[4] ;
  wire \r9_reg_n_0_[5] ;
  wire \r9_reg_n_0_[6] ;
  wire \r9_reg_n_0_[7] ;
  wire \r9_reg_n_0_[8] ;
  wire \r9_reg_n_0_[9] ;

  IBUF \A1_IBUF[0]_inst 
       (.I(A1[0]),
        .O(A1_IBUF[0]));
  IBUF \A1_IBUF[1]_inst 
       (.I(A1[1]),
        .O(A1_IBUF[1]));
  IBUF \A1_IBUF[2]_inst 
       (.I(A1[2]),
        .O(A1_IBUF[2]));
  IBUF \A1_IBUF[3]_inst 
       (.I(A1[3]),
        .O(A1_IBUF[3]));
  IBUF \A1_IBUF[4]_inst 
       (.I(A1[4]),
        .O(A1_IBUF[4]));
  IBUF \A2_IBUF[0]_inst 
       (.I(A2[0]),
        .O(A2_IBUF[0]));
  IBUF \A2_IBUF[1]_inst 
       (.I(A2[1]),
        .O(A2_IBUF[1]));
  IBUF \A2_IBUF[2]_inst 
       (.I(A2[2]),
        .O(A2_IBUF[2]));
  IBUF \A2_IBUF[3]_inst 
       (.I(A2[3]),
        .O(A2_IBUF[3]));
  IBUF \A2_IBUF[4]_inst 
       (.I(A2[4]),
        .O(A2_IBUF[4]));
  IBUF \A3_IBUF[0]_inst 
       (.I(A3[0]),
        .O(A3_IBUF[0]));
  IBUF \A3_IBUF[1]_inst 
       (.I(A3[1]),
        .O(A3_IBUF[1]));
  IBUF \A3_IBUF[2]_inst 
       (.I(A3[2]),
        .O(A3_IBUF[2]));
  IBUF \A3_IBUF[3]_inst 
       (.I(A3[3]),
        .O(A3_IBUF[3]));
  IBUF \A3_IBUF[4]_inst 
       (.I(A3[4]),
        .O(A3_IBUF[4]));
  GND GND
       (.G(\<const0> ));
  OBUF \RD1_OBUF[0]_inst 
       (.I(RD1_OBUF[0]),
        .O(RD1[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_1 
       (.I0(\RD1_OBUF[0]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[0]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[0]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[0]_inst_i_5_n_0 ),
        .O(RD1_OBUF[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_10 
       (.I0(\r11_reg_n_0_[0] ),
        .I1(\r10_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_11 
       (.I0(\r15_reg_n_0_[0] ),
        .I1(\r14_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[0]_inst_i_12 
       (.I0(\r3_reg_n_0_[0] ),
        .I1(\r2_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_13 
       (.I0(\r7_reg_n_0_[0] ),
        .I1(\r6_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[0]_inst_i_2 
       (.I0(\RD1_OBUF[0]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[0]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[0]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[0]_inst_i_3 
       (.I0(\RD1_OBUF[0]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[0]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[0]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[0]_inst_i_4 
       (.I0(\RD1_OBUF[0]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[0]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[0]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[0]_inst_i_5 
       (.I0(\RD1_OBUF[0]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[0]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[0]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_6 
       (.I0(\r27_reg_n_0_[0] ),
        .I1(\r26_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_7 
       (.I0(\r31_reg_n_0_[0] ),
        .I1(\r30_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_8 
       (.I0(\r19_reg_n_0_[0] ),
        .I1(\r18_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[0]_inst_i_9 
       (.I0(\r23_reg_n_0_[0] ),
        .I1(\r22_reg_n_0_[0] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[0] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[0] ),
        .O(\RD1_OBUF[0]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[10]_inst 
       (.I(RD1_OBUF[10]),
        .O(RD1[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_1 
       (.I0(\RD1_OBUF[10]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[10]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[10]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[10]_inst_i_5_n_0 ),
        .O(RD1_OBUF[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_10 
       (.I0(\r11_reg_n_0_[10] ),
        .I1(\r10_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_11 
       (.I0(\r15_reg_n_0_[10] ),
        .I1(\r14_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[10]_inst_i_12 
       (.I0(\r3_reg_n_0_[10] ),
        .I1(\r2_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_13 
       (.I0(\r7_reg_n_0_[10] ),
        .I1(\r6_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[10]_inst_i_2 
       (.I0(\RD1_OBUF[10]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[10]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[10]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[10]_inst_i_3 
       (.I0(\RD1_OBUF[10]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[10]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[10]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[10]_inst_i_4 
       (.I0(\RD1_OBUF[10]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[10]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[10]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[10]_inst_i_5 
       (.I0(\RD1_OBUF[10]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[10]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[10]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_6 
       (.I0(\r27_reg_n_0_[10] ),
        .I1(\r26_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_7 
       (.I0(\r31_reg_n_0_[10] ),
        .I1(\r30_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_8 
       (.I0(\r19_reg_n_0_[10] ),
        .I1(\r18_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[10]_inst_i_9 
       (.I0(\r23_reg_n_0_[10] ),
        .I1(\r22_reg_n_0_[10] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[10] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[10] ),
        .O(\RD1_OBUF[10]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[11]_inst 
       (.I(RD1_OBUF[11]),
        .O(RD1[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_1 
       (.I0(\RD1_OBUF[11]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[11]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[11]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[11]_inst_i_5_n_0 ),
        .O(RD1_OBUF[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_10 
       (.I0(\r11_reg_n_0_[11] ),
        .I1(\r10_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_11 
       (.I0(\r15_reg_n_0_[11] ),
        .I1(\r14_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[11]_inst_i_12 
       (.I0(\r3_reg_n_0_[11] ),
        .I1(\r2_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_13 
       (.I0(\r7_reg_n_0_[11] ),
        .I1(\r6_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[11]_inst_i_2 
       (.I0(\RD1_OBUF[11]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[11]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[11]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[11]_inst_i_3 
       (.I0(\RD1_OBUF[11]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[11]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[11]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[11]_inst_i_4 
       (.I0(\RD1_OBUF[11]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[11]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[11]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[11]_inst_i_5 
       (.I0(\RD1_OBUF[11]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[11]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[11]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_6 
       (.I0(\r27_reg_n_0_[11] ),
        .I1(\r26_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_7 
       (.I0(\r31_reg_n_0_[11] ),
        .I1(\r30_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_8 
       (.I0(\r19_reg_n_0_[11] ),
        .I1(\r18_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[11]_inst_i_9 
       (.I0(\r23_reg_n_0_[11] ),
        .I1(\r22_reg_n_0_[11] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[11] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[11] ),
        .O(\RD1_OBUF[11]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[12]_inst 
       (.I(RD1_OBUF[12]),
        .O(RD1[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_1 
       (.I0(\RD1_OBUF[12]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[12]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[12]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[12]_inst_i_5_n_0 ),
        .O(RD1_OBUF[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_10 
       (.I0(\r11_reg_n_0_[12] ),
        .I1(\r10_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_11 
       (.I0(\r15_reg_n_0_[12] ),
        .I1(\r14_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[12]_inst_i_12 
       (.I0(\r3_reg_n_0_[12] ),
        .I1(\r2_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_13 
       (.I0(\r7_reg_n_0_[12] ),
        .I1(\r6_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[12]_inst_i_2 
       (.I0(\RD1_OBUF[12]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[12]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[12]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[12]_inst_i_3 
       (.I0(\RD1_OBUF[12]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[12]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[12]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[12]_inst_i_4 
       (.I0(\RD1_OBUF[12]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[12]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[12]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[12]_inst_i_5 
       (.I0(\RD1_OBUF[12]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[12]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[12]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_6 
       (.I0(\r27_reg_n_0_[12] ),
        .I1(\r26_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_7 
       (.I0(\r31_reg_n_0_[12] ),
        .I1(\r30_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_8 
       (.I0(\r19_reg_n_0_[12] ),
        .I1(\r18_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[12]_inst_i_9 
       (.I0(\r23_reg_n_0_[12] ),
        .I1(\r22_reg_n_0_[12] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[12] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[12] ),
        .O(\RD1_OBUF[12]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[13]_inst 
       (.I(RD1_OBUF[13]),
        .O(RD1[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_1 
       (.I0(\RD1_OBUF[13]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[13]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[13]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[13]_inst_i_5_n_0 ),
        .O(RD1_OBUF[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_10 
       (.I0(\r11_reg_n_0_[13] ),
        .I1(\r10_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_11 
       (.I0(\r15_reg_n_0_[13] ),
        .I1(\r14_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[13]_inst_i_12 
       (.I0(\r3_reg_n_0_[13] ),
        .I1(\r2_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_13 
       (.I0(\r7_reg_n_0_[13] ),
        .I1(\r6_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[13]_inst_i_2 
       (.I0(\RD1_OBUF[13]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[13]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[13]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[13]_inst_i_3 
       (.I0(\RD1_OBUF[13]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[13]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[13]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[13]_inst_i_4 
       (.I0(\RD1_OBUF[13]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[13]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[13]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[13]_inst_i_5 
       (.I0(\RD1_OBUF[13]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[13]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[13]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_6 
       (.I0(\r27_reg_n_0_[13] ),
        .I1(\r26_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_7 
       (.I0(\r31_reg_n_0_[13] ),
        .I1(\r30_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_8 
       (.I0(\r19_reg_n_0_[13] ),
        .I1(\r18_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[13]_inst_i_9 
       (.I0(\r23_reg_n_0_[13] ),
        .I1(\r22_reg_n_0_[13] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[13] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[13] ),
        .O(\RD1_OBUF[13]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[14]_inst 
       (.I(RD1_OBUF[14]),
        .O(RD1[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_1 
       (.I0(\RD1_OBUF[14]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[14]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[14]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[14]_inst_i_5_n_0 ),
        .O(RD1_OBUF[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_10 
       (.I0(\r11_reg_n_0_[14] ),
        .I1(\r10_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_11 
       (.I0(\r15_reg_n_0_[14] ),
        .I1(\r14_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[14]_inst_i_12 
       (.I0(\r3_reg_n_0_[14] ),
        .I1(\r2_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_13 
       (.I0(\r7_reg_n_0_[14] ),
        .I1(\r6_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[14]_inst_i_2 
       (.I0(\RD1_OBUF[14]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[14]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[14]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[14]_inst_i_3 
       (.I0(\RD1_OBUF[14]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[14]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[14]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[14]_inst_i_4 
       (.I0(\RD1_OBUF[14]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[14]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[14]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[14]_inst_i_5 
       (.I0(\RD1_OBUF[14]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[14]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[14]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_6 
       (.I0(\r27_reg_n_0_[14] ),
        .I1(\r26_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_7 
       (.I0(\r31_reg_n_0_[14] ),
        .I1(\r30_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_8 
       (.I0(\r19_reg_n_0_[14] ),
        .I1(\r18_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[14]_inst_i_9 
       (.I0(\r23_reg_n_0_[14] ),
        .I1(\r22_reg_n_0_[14] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[14] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[14] ),
        .O(\RD1_OBUF[14]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[15]_inst 
       (.I(RD1_OBUF[15]),
        .O(RD1[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_1 
       (.I0(\RD1_OBUF[15]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[15]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[15]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[15]_inst_i_5_n_0 ),
        .O(RD1_OBUF[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_10 
       (.I0(\r11_reg_n_0_[15] ),
        .I1(\r10_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_11 
       (.I0(\r15_reg_n_0_[15] ),
        .I1(\r14_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[15]_inst_i_12 
       (.I0(\r3_reg_n_0_[15] ),
        .I1(\r2_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_13 
       (.I0(\r7_reg_n_0_[15] ),
        .I1(\r6_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[15]_inst_i_2 
       (.I0(\RD1_OBUF[15]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[15]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[15]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[15]_inst_i_3 
       (.I0(\RD1_OBUF[15]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[15]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[15]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[15]_inst_i_4 
       (.I0(\RD1_OBUF[15]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[15]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[15]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[15]_inst_i_5 
       (.I0(\RD1_OBUF[15]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[15]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[15]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_6 
       (.I0(\r27_reg_n_0_[15] ),
        .I1(\r26_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_7 
       (.I0(\r31_reg_n_0_[15] ),
        .I1(\r30_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_8 
       (.I0(\r19_reg_n_0_[15] ),
        .I1(\r18_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[15]_inst_i_9 
       (.I0(\r23_reg_n_0_[15] ),
        .I1(\r22_reg_n_0_[15] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[15] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[15] ),
        .O(\RD1_OBUF[15]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[16]_inst 
       (.I(RD1_OBUF[16]),
        .O(RD1[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_1 
       (.I0(\RD1_OBUF[16]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[16]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[16]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[16]_inst_i_5_n_0 ),
        .O(RD1_OBUF[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_10 
       (.I0(\r11_reg_n_0_[16] ),
        .I1(\r10_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_11 
       (.I0(\r15_reg_n_0_[16] ),
        .I1(\r14_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[16]_inst_i_12 
       (.I0(\r3_reg_n_0_[16] ),
        .I1(\r2_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_13 
       (.I0(\r7_reg_n_0_[16] ),
        .I1(\r6_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[16]_inst_i_2 
       (.I0(\RD1_OBUF[16]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[16]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[16]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[16]_inst_i_3 
       (.I0(\RD1_OBUF[16]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[16]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[16]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[16]_inst_i_4 
       (.I0(\RD1_OBUF[16]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[16]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[16]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[16]_inst_i_5 
       (.I0(\RD1_OBUF[16]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[16]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[16]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_6 
       (.I0(\r27_reg_n_0_[16] ),
        .I1(\r26_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_7 
       (.I0(\r31_reg_n_0_[16] ),
        .I1(\r30_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_8 
       (.I0(\r19_reg_n_0_[16] ),
        .I1(\r18_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[16]_inst_i_9 
       (.I0(\r23_reg_n_0_[16] ),
        .I1(\r22_reg_n_0_[16] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[16] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[16] ),
        .O(\RD1_OBUF[16]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[17]_inst 
       (.I(RD1_OBUF[17]),
        .O(RD1[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_1 
       (.I0(\RD1_OBUF[17]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[17]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[17]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[17]_inst_i_5_n_0 ),
        .O(RD1_OBUF[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_10 
       (.I0(\r11_reg_n_0_[17] ),
        .I1(\r10_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_11 
       (.I0(\r15_reg_n_0_[17] ),
        .I1(\r14_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[17]_inst_i_12 
       (.I0(\r3_reg_n_0_[17] ),
        .I1(\r2_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_13 
       (.I0(\r7_reg_n_0_[17] ),
        .I1(\r6_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[17]_inst_i_2 
       (.I0(\RD1_OBUF[17]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[17]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[17]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[17]_inst_i_3 
       (.I0(\RD1_OBUF[17]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[17]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[17]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[17]_inst_i_4 
       (.I0(\RD1_OBUF[17]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[17]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[17]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[17]_inst_i_5 
       (.I0(\RD1_OBUF[17]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[17]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[17]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_6 
       (.I0(\r27_reg_n_0_[17] ),
        .I1(\r26_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_7 
       (.I0(\r31_reg_n_0_[17] ),
        .I1(\r30_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_8 
       (.I0(\r19_reg_n_0_[17] ),
        .I1(\r18_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[17]_inst_i_9 
       (.I0(\r23_reg_n_0_[17] ),
        .I1(\r22_reg_n_0_[17] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[17] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[17] ),
        .O(\RD1_OBUF[17]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[18]_inst 
       (.I(RD1_OBUF[18]),
        .O(RD1[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_1 
       (.I0(\RD1_OBUF[18]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[18]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[18]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[18]_inst_i_5_n_0 ),
        .O(RD1_OBUF[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_10 
       (.I0(\r11_reg_n_0_[18] ),
        .I1(\r10_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_11 
       (.I0(\r15_reg_n_0_[18] ),
        .I1(\r14_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[18]_inst_i_12 
       (.I0(\r3_reg_n_0_[18] ),
        .I1(\r2_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_13 
       (.I0(\r7_reg_n_0_[18] ),
        .I1(\r6_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[18]_inst_i_2 
       (.I0(\RD1_OBUF[18]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[18]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[18]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[18]_inst_i_3 
       (.I0(\RD1_OBUF[18]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[18]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[18]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[18]_inst_i_4 
       (.I0(\RD1_OBUF[18]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[18]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[18]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[18]_inst_i_5 
       (.I0(\RD1_OBUF[18]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[18]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[18]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_6 
       (.I0(\r27_reg_n_0_[18] ),
        .I1(\r26_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_7 
       (.I0(\r31_reg_n_0_[18] ),
        .I1(\r30_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_8 
       (.I0(\r19_reg_n_0_[18] ),
        .I1(\r18_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[18]_inst_i_9 
       (.I0(\r23_reg_n_0_[18] ),
        .I1(\r22_reg_n_0_[18] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[18] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[18] ),
        .O(\RD1_OBUF[18]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[19]_inst 
       (.I(RD1_OBUF[19]),
        .O(RD1[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_1 
       (.I0(\RD1_OBUF[19]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[19]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[19]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[19]_inst_i_5_n_0 ),
        .O(RD1_OBUF[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_10 
       (.I0(\r11_reg_n_0_[19] ),
        .I1(\r10_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_11 
       (.I0(\r15_reg_n_0_[19] ),
        .I1(\r14_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[19]_inst_i_12 
       (.I0(\r3_reg_n_0_[19] ),
        .I1(\r2_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_13 
       (.I0(\r7_reg_n_0_[19] ),
        .I1(\r6_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[19]_inst_i_2 
       (.I0(\RD1_OBUF[19]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[19]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[19]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[19]_inst_i_3 
       (.I0(\RD1_OBUF[19]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[19]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[19]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[19]_inst_i_4 
       (.I0(\RD1_OBUF[19]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[19]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[19]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[19]_inst_i_5 
       (.I0(\RD1_OBUF[19]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[19]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[19]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_6 
       (.I0(\r27_reg_n_0_[19] ),
        .I1(\r26_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_7 
       (.I0(\r31_reg_n_0_[19] ),
        .I1(\r30_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_8 
       (.I0(\r19_reg_n_0_[19] ),
        .I1(\r18_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[19]_inst_i_9 
       (.I0(\r23_reg_n_0_[19] ),
        .I1(\r22_reg_n_0_[19] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[19] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[19] ),
        .O(\RD1_OBUF[19]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[1]_inst 
       (.I(RD1_OBUF[1]),
        .O(RD1[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_1 
       (.I0(\RD1_OBUF[1]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[1]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[1]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[1]_inst_i_5_n_0 ),
        .O(RD1_OBUF[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_10 
       (.I0(\r11_reg_n_0_[1] ),
        .I1(\r10_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_11 
       (.I0(\r15_reg_n_0_[1] ),
        .I1(\r14_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[1]_inst_i_12 
       (.I0(\r3_reg_n_0_[1] ),
        .I1(\r2_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_13 
       (.I0(\r7_reg_n_0_[1] ),
        .I1(\r6_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[1]_inst_i_2 
       (.I0(\RD1_OBUF[1]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[1]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[1]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[1]_inst_i_3 
       (.I0(\RD1_OBUF[1]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[1]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[1]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[1]_inst_i_4 
       (.I0(\RD1_OBUF[1]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[1]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[1]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[1]_inst_i_5 
       (.I0(\RD1_OBUF[1]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[1]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[1]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_6 
       (.I0(\r27_reg_n_0_[1] ),
        .I1(\r26_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_7 
       (.I0(\r31_reg_n_0_[1] ),
        .I1(\r30_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_8 
       (.I0(\r19_reg_n_0_[1] ),
        .I1(\r18_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[1]_inst_i_9 
       (.I0(\r23_reg_n_0_[1] ),
        .I1(\r22_reg_n_0_[1] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[1] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[1] ),
        .O(\RD1_OBUF[1]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[20]_inst 
       (.I(RD1_OBUF[20]),
        .O(RD1[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_1 
       (.I0(\RD1_OBUF[20]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[20]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[20]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[20]_inst_i_5_n_0 ),
        .O(RD1_OBUF[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_10 
       (.I0(\r11_reg_n_0_[20] ),
        .I1(\r10_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_11 
       (.I0(\r15_reg_n_0_[20] ),
        .I1(\r14_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[20]_inst_i_12 
       (.I0(\r3_reg_n_0_[20] ),
        .I1(\r2_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_13 
       (.I0(\r7_reg_n_0_[20] ),
        .I1(\r6_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[20]_inst_i_2 
       (.I0(\RD1_OBUF[20]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[20]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[20]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[20]_inst_i_3 
       (.I0(\RD1_OBUF[20]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[20]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[20]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[20]_inst_i_4 
       (.I0(\RD1_OBUF[20]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[20]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[20]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[20]_inst_i_5 
       (.I0(\RD1_OBUF[20]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[20]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[20]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_6 
       (.I0(\r27_reg_n_0_[20] ),
        .I1(\r26_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_7 
       (.I0(\r31_reg_n_0_[20] ),
        .I1(\r30_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_8 
       (.I0(\r19_reg_n_0_[20] ),
        .I1(\r18_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[20]_inst_i_9 
       (.I0(\r23_reg_n_0_[20] ),
        .I1(\r22_reg_n_0_[20] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[20] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[20] ),
        .O(\RD1_OBUF[20]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[21]_inst 
       (.I(RD1_OBUF[21]),
        .O(RD1[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_1 
       (.I0(\RD1_OBUF[21]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[21]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[21]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[21]_inst_i_5_n_0 ),
        .O(RD1_OBUF[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_10 
       (.I0(\r11_reg_n_0_[21] ),
        .I1(\r10_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_11 
       (.I0(\r15_reg_n_0_[21] ),
        .I1(\r14_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[21]_inst_i_12 
       (.I0(\r3_reg_n_0_[21] ),
        .I1(\r2_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_13 
       (.I0(\r7_reg_n_0_[21] ),
        .I1(\r6_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[21]_inst_i_2 
       (.I0(\RD1_OBUF[21]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[21]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[21]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[21]_inst_i_3 
       (.I0(\RD1_OBUF[21]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[21]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[21]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[21]_inst_i_4 
       (.I0(\RD1_OBUF[21]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[21]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[21]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[21]_inst_i_5 
       (.I0(\RD1_OBUF[21]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[21]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[21]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_6 
       (.I0(\r27_reg_n_0_[21] ),
        .I1(\r26_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_7 
       (.I0(\r31_reg_n_0_[21] ),
        .I1(\r30_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_8 
       (.I0(\r19_reg_n_0_[21] ),
        .I1(\r18_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[21]_inst_i_9 
       (.I0(\r23_reg_n_0_[21] ),
        .I1(\r22_reg_n_0_[21] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[21] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[21] ),
        .O(\RD1_OBUF[21]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[22]_inst 
       (.I(RD1_OBUF[22]),
        .O(RD1[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_1 
       (.I0(\RD1_OBUF[22]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[22]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[22]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[22]_inst_i_5_n_0 ),
        .O(RD1_OBUF[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_10 
       (.I0(\r11_reg_n_0_[22] ),
        .I1(\r10_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_11 
       (.I0(\r15_reg_n_0_[22] ),
        .I1(\r14_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[22]_inst_i_12 
       (.I0(\r3_reg_n_0_[22] ),
        .I1(\r2_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_13 
       (.I0(\r7_reg_n_0_[22] ),
        .I1(\r6_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[22]_inst_i_2 
       (.I0(\RD1_OBUF[22]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[22]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[22]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[22]_inst_i_3 
       (.I0(\RD1_OBUF[22]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[22]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[22]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[22]_inst_i_4 
       (.I0(\RD1_OBUF[22]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[22]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[22]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[22]_inst_i_5 
       (.I0(\RD1_OBUF[22]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[22]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[22]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_6 
       (.I0(\r27_reg_n_0_[22] ),
        .I1(\r26_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_7 
       (.I0(\r31_reg_n_0_[22] ),
        .I1(\r30_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_8 
       (.I0(\r19_reg_n_0_[22] ),
        .I1(\r18_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[22]_inst_i_9 
       (.I0(\r23_reg_n_0_[22] ),
        .I1(\r22_reg_n_0_[22] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[22] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[22] ),
        .O(\RD1_OBUF[22]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[23]_inst 
       (.I(RD1_OBUF[23]),
        .O(RD1[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_1 
       (.I0(\RD1_OBUF[23]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[23]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[23]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[23]_inst_i_5_n_0 ),
        .O(RD1_OBUF[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_10 
       (.I0(\r11_reg_n_0_[23] ),
        .I1(\r10_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_11 
       (.I0(\r15_reg_n_0_[23] ),
        .I1(\r14_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[23]_inst_i_12 
       (.I0(\r3_reg_n_0_[23] ),
        .I1(\r2_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_13 
       (.I0(\r7_reg_n_0_[23] ),
        .I1(\r6_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[23]_inst_i_2 
       (.I0(\RD1_OBUF[23]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[23]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[23]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[23]_inst_i_3 
       (.I0(\RD1_OBUF[23]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[23]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[23]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[23]_inst_i_4 
       (.I0(\RD1_OBUF[23]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[23]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[23]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[23]_inst_i_5 
       (.I0(\RD1_OBUF[23]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[23]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[23]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_6 
       (.I0(\r27_reg_n_0_[23] ),
        .I1(\r26_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_7 
       (.I0(\r31_reg_n_0_[23] ),
        .I1(\r30_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_8 
       (.I0(\r19_reg_n_0_[23] ),
        .I1(\r18_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[23]_inst_i_9 
       (.I0(\r23_reg_n_0_[23] ),
        .I1(\r22_reg_n_0_[23] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[23] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[23] ),
        .O(\RD1_OBUF[23]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[24]_inst 
       (.I(RD1_OBUF[24]),
        .O(RD1[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_1 
       (.I0(\RD1_OBUF[24]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[24]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[24]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[24]_inst_i_5_n_0 ),
        .O(RD1_OBUF[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_10 
       (.I0(\r11_reg_n_0_[24] ),
        .I1(\r10_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_11 
       (.I0(\r15_reg_n_0_[24] ),
        .I1(\r14_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[24]_inst_i_12 
       (.I0(\r3_reg_n_0_[24] ),
        .I1(\r2_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_13 
       (.I0(\r7_reg_n_0_[24] ),
        .I1(\r6_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[24]_inst_i_2 
       (.I0(\RD1_OBUF[24]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[24]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[24]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[24]_inst_i_3 
       (.I0(\RD1_OBUF[24]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[24]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[24]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[24]_inst_i_4 
       (.I0(\RD1_OBUF[24]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[24]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[24]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[24]_inst_i_5 
       (.I0(\RD1_OBUF[24]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[24]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[24]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_6 
       (.I0(\r27_reg_n_0_[24] ),
        .I1(\r26_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_7 
       (.I0(\r31_reg_n_0_[24] ),
        .I1(\r30_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_8 
       (.I0(\r19_reg_n_0_[24] ),
        .I1(\r18_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[24]_inst_i_9 
       (.I0(\r23_reg_n_0_[24] ),
        .I1(\r22_reg_n_0_[24] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[24] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[24] ),
        .O(\RD1_OBUF[24]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[25]_inst 
       (.I(RD1_OBUF[25]),
        .O(RD1[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_1 
       (.I0(\RD1_OBUF[25]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[25]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[25]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[25]_inst_i_5_n_0 ),
        .O(RD1_OBUF[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_10 
       (.I0(\r11_reg_n_0_[25] ),
        .I1(\r10_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_11 
       (.I0(\r15_reg_n_0_[25] ),
        .I1(\r14_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[25]_inst_i_12 
       (.I0(\r3_reg_n_0_[25] ),
        .I1(\r2_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_13 
       (.I0(\r7_reg_n_0_[25] ),
        .I1(\r6_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[25]_inst_i_2 
       (.I0(\RD1_OBUF[25]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[25]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[25]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[25]_inst_i_3 
       (.I0(\RD1_OBUF[25]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[25]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[25]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[25]_inst_i_4 
       (.I0(\RD1_OBUF[25]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[25]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[25]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[25]_inst_i_5 
       (.I0(\RD1_OBUF[25]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[25]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[25]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_6 
       (.I0(\r27_reg_n_0_[25] ),
        .I1(\r26_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_7 
       (.I0(\r31_reg_n_0_[25] ),
        .I1(\r30_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_8 
       (.I0(\r19_reg_n_0_[25] ),
        .I1(\r18_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[25]_inst_i_9 
       (.I0(\r23_reg_n_0_[25] ),
        .I1(\r22_reg_n_0_[25] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[25] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[25] ),
        .O(\RD1_OBUF[25]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[26]_inst 
       (.I(RD1_OBUF[26]),
        .O(RD1[26]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_1 
       (.I0(\RD1_OBUF[26]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[26]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[26]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[26]_inst_i_5_n_0 ),
        .O(RD1_OBUF[26]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_10 
       (.I0(\r11_reg_n_0_[26] ),
        .I1(\r10_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_11 
       (.I0(\r15_reg_n_0_[26] ),
        .I1(\r14_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[26]_inst_i_12 
       (.I0(\r3_reg_n_0_[26] ),
        .I1(\r2_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_13 
       (.I0(\r7_reg_n_0_[26] ),
        .I1(\r6_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[26]_inst_i_2 
       (.I0(\RD1_OBUF[26]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[26]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[26]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[26]_inst_i_3 
       (.I0(\RD1_OBUF[26]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[26]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[26]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[26]_inst_i_4 
       (.I0(\RD1_OBUF[26]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[26]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[26]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[26]_inst_i_5 
       (.I0(\RD1_OBUF[26]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[26]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[26]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_6 
       (.I0(\r27_reg_n_0_[26] ),
        .I1(\r26_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_7 
       (.I0(\r31_reg_n_0_[26] ),
        .I1(\r30_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_8 
       (.I0(\r19_reg_n_0_[26] ),
        .I1(\r18_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[26]_inst_i_9 
       (.I0(\r23_reg_n_0_[26] ),
        .I1(\r22_reg_n_0_[26] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[26] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[26] ),
        .O(\RD1_OBUF[26]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[27]_inst 
       (.I(RD1_OBUF[27]),
        .O(RD1[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_1 
       (.I0(\RD1_OBUF[27]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[27]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[27]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[27]_inst_i_5_n_0 ),
        .O(RD1_OBUF[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_10 
       (.I0(\r11_reg_n_0_[27] ),
        .I1(\r10_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_11 
       (.I0(\r15_reg_n_0_[27] ),
        .I1(\r14_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[27]_inst_i_12 
       (.I0(\r3_reg_n_0_[27] ),
        .I1(\r2_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_13 
       (.I0(\r7_reg_n_0_[27] ),
        .I1(\r6_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[27]_inst_i_2 
       (.I0(\RD1_OBUF[27]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[27]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[27]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[27]_inst_i_3 
       (.I0(\RD1_OBUF[27]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[27]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[27]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[27]_inst_i_4 
       (.I0(\RD1_OBUF[27]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[27]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[27]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[27]_inst_i_5 
       (.I0(\RD1_OBUF[27]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[27]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[27]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_6 
       (.I0(\r27_reg_n_0_[27] ),
        .I1(\r26_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_7 
       (.I0(\r31_reg_n_0_[27] ),
        .I1(\r30_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_8 
       (.I0(\r19_reg_n_0_[27] ),
        .I1(\r18_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[27]_inst_i_9 
       (.I0(\r23_reg_n_0_[27] ),
        .I1(\r22_reg_n_0_[27] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[27] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[27] ),
        .O(\RD1_OBUF[27]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[28]_inst 
       (.I(RD1_OBUF[28]),
        .O(RD1[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_1 
       (.I0(\RD1_OBUF[28]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[28]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[28]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[28]_inst_i_5_n_0 ),
        .O(RD1_OBUF[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_10 
       (.I0(\r11_reg_n_0_[28] ),
        .I1(\r10_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_11 
       (.I0(\r15_reg_n_0_[28] ),
        .I1(\r14_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[28]_inst_i_12 
       (.I0(\r3_reg_n_0_[28] ),
        .I1(\r2_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_13 
       (.I0(\r7_reg_n_0_[28] ),
        .I1(\r6_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[28]_inst_i_2 
       (.I0(\RD1_OBUF[28]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[28]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[28]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[28]_inst_i_3 
       (.I0(\RD1_OBUF[28]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[28]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[28]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[28]_inst_i_4 
       (.I0(\RD1_OBUF[28]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[28]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[28]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[28]_inst_i_5 
       (.I0(\RD1_OBUF[28]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[28]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[28]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_6 
       (.I0(\r27_reg_n_0_[28] ),
        .I1(\r26_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_7 
       (.I0(\r31_reg_n_0_[28] ),
        .I1(\r30_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_8 
       (.I0(\r19_reg_n_0_[28] ),
        .I1(\r18_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[28]_inst_i_9 
       (.I0(\r23_reg_n_0_[28] ),
        .I1(\r22_reg_n_0_[28] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[28] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[28] ),
        .O(\RD1_OBUF[28]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[29]_inst 
       (.I(RD1_OBUF[29]),
        .O(RD1[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_1 
       (.I0(\RD1_OBUF[29]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[29]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[29]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[29]_inst_i_5_n_0 ),
        .O(RD1_OBUF[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_10 
       (.I0(\r11_reg_n_0_[29] ),
        .I1(\r10_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_11 
       (.I0(\r15_reg_n_0_[29] ),
        .I1(\r14_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[29]_inst_i_12 
       (.I0(\r3_reg_n_0_[29] ),
        .I1(\r2_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_13 
       (.I0(\r7_reg_n_0_[29] ),
        .I1(\r6_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[29]_inst_i_2 
       (.I0(\RD1_OBUF[29]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[29]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[29]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[29]_inst_i_3 
       (.I0(\RD1_OBUF[29]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[29]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[29]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[29]_inst_i_4 
       (.I0(\RD1_OBUF[29]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[29]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[29]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[29]_inst_i_5 
       (.I0(\RD1_OBUF[29]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[29]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[29]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_6 
       (.I0(\r27_reg_n_0_[29] ),
        .I1(\r26_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_7 
       (.I0(\r31_reg_n_0_[29] ),
        .I1(\r30_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_8 
       (.I0(\r19_reg_n_0_[29] ),
        .I1(\r18_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[29]_inst_i_9 
       (.I0(\r23_reg_n_0_[29] ),
        .I1(\r22_reg_n_0_[29] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[29] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[29] ),
        .O(\RD1_OBUF[29]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[2]_inst 
       (.I(RD1_OBUF[2]),
        .O(RD1[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_1 
       (.I0(\RD1_OBUF[2]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[2]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[2]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[2]_inst_i_5_n_0 ),
        .O(RD1_OBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_10 
       (.I0(\r11_reg_n_0_[2] ),
        .I1(\r10_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_11 
       (.I0(\r15_reg_n_0_[2] ),
        .I1(\r14_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[2]_inst_i_12 
       (.I0(\r3_reg_n_0_[2] ),
        .I1(\r2_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_13 
       (.I0(\r7_reg_n_0_[2] ),
        .I1(\r6_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[2]_inst_i_2 
       (.I0(\RD1_OBUF[2]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[2]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[2]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[2]_inst_i_3 
       (.I0(\RD1_OBUF[2]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[2]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[2]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[2]_inst_i_4 
       (.I0(\RD1_OBUF[2]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[2]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[2]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[2]_inst_i_5 
       (.I0(\RD1_OBUF[2]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[2]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[2]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_6 
       (.I0(\r27_reg_n_0_[2] ),
        .I1(\r26_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_7 
       (.I0(\r31_reg_n_0_[2] ),
        .I1(\r30_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_8 
       (.I0(\r19_reg_n_0_[2] ),
        .I1(\r18_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[2]_inst_i_9 
       (.I0(\r23_reg_n_0_[2] ),
        .I1(\r22_reg_n_0_[2] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[2] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[2] ),
        .O(\RD1_OBUF[2]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[30]_inst 
       (.I(RD1_OBUF[30]),
        .O(RD1[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_1 
       (.I0(\RD1_OBUF[30]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[30]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[30]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[30]_inst_i_5_n_0 ),
        .O(RD1_OBUF[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_10 
       (.I0(\r11_reg_n_0_[30] ),
        .I1(\r10_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_11 
       (.I0(\r15_reg_n_0_[30] ),
        .I1(\r14_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[30]_inst_i_12 
       (.I0(\r3_reg_n_0_[30] ),
        .I1(\r2_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_13 
       (.I0(\r7_reg_n_0_[30] ),
        .I1(\r6_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[30]_inst_i_2 
       (.I0(\RD1_OBUF[30]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[30]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[30]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[30]_inst_i_3 
       (.I0(\RD1_OBUF[30]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[30]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[30]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[30]_inst_i_4 
       (.I0(\RD1_OBUF[30]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[30]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[30]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[30]_inst_i_5 
       (.I0(\RD1_OBUF[30]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[30]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[30]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_6 
       (.I0(\r27_reg_n_0_[30] ),
        .I1(\r26_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_7 
       (.I0(\r31_reg_n_0_[30] ),
        .I1(\r30_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_8 
       (.I0(\r19_reg_n_0_[30] ),
        .I1(\r18_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[30]_inst_i_9 
       (.I0(\r23_reg_n_0_[30] ),
        .I1(\r22_reg_n_0_[30] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[30] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[30] ),
        .O(\RD1_OBUF[30]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[31]_inst 
       (.I(RD1_OBUF[31]),
        .O(RD1[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_1 
       (.I0(\RD1_OBUF[31]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[31]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[31]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[31]_inst_i_5_n_0 ),
        .O(RD1_OBUF[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_10 
       (.I0(\r11_reg_n_0_[31] ),
        .I1(\r10_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_11 
       (.I0(\r15_reg_n_0_[31] ),
        .I1(\r14_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[31]_inst_i_12 
       (.I0(\r3_reg_n_0_[31] ),
        .I1(\r2_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_13 
       (.I0(\r7_reg_n_0_[31] ),
        .I1(\r6_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[31]_inst_i_2 
       (.I0(\RD1_OBUF[31]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[31]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[31]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[31]_inst_i_3 
       (.I0(\RD1_OBUF[31]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[31]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[31]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[31]_inst_i_4 
       (.I0(\RD1_OBUF[31]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[31]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[31]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[31]_inst_i_5 
       (.I0(\RD1_OBUF[31]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[31]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[31]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_6 
       (.I0(\r27_reg_n_0_[31] ),
        .I1(\r26_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_7 
       (.I0(\r31_reg_n_0_[31] ),
        .I1(\r30_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_8 
       (.I0(\r19_reg_n_0_[31] ),
        .I1(\r18_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[31]_inst_i_9 
       (.I0(\r23_reg_n_0_[31] ),
        .I1(\r22_reg_n_0_[31] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[31] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[31] ),
        .O(\RD1_OBUF[31]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[3]_inst 
       (.I(RD1_OBUF[3]),
        .O(RD1[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_1 
       (.I0(\RD1_OBUF[3]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[3]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[3]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[3]_inst_i_5_n_0 ),
        .O(RD1_OBUF[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_10 
       (.I0(\r11_reg_n_0_[3] ),
        .I1(\r10_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_11 
       (.I0(\r15_reg_n_0_[3] ),
        .I1(\r14_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[3]_inst_i_12 
       (.I0(\r3_reg_n_0_[3] ),
        .I1(\r2_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_13 
       (.I0(\r7_reg_n_0_[3] ),
        .I1(\r6_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[3]_inst_i_2 
       (.I0(\RD1_OBUF[3]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[3]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[3]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[3]_inst_i_3 
       (.I0(\RD1_OBUF[3]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[3]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[3]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[3]_inst_i_4 
       (.I0(\RD1_OBUF[3]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[3]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[3]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[3]_inst_i_5 
       (.I0(\RD1_OBUF[3]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[3]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[3]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_6 
       (.I0(\r27_reg_n_0_[3] ),
        .I1(\r26_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_7 
       (.I0(\r31_reg_n_0_[3] ),
        .I1(\r30_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_8 
       (.I0(\r19_reg_n_0_[3] ),
        .I1(\r18_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[3]_inst_i_9 
       (.I0(\r23_reg_n_0_[3] ),
        .I1(\r22_reg_n_0_[3] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[3] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[3] ),
        .O(\RD1_OBUF[3]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[4]_inst 
       (.I(RD1_OBUF[4]),
        .O(RD1[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_1 
       (.I0(\RD1_OBUF[4]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[4]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[4]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[4]_inst_i_5_n_0 ),
        .O(RD1_OBUF[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_10 
       (.I0(\r11_reg_n_0_[4] ),
        .I1(\r10_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_11 
       (.I0(\r15_reg_n_0_[4] ),
        .I1(\r14_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[4]_inst_i_12 
       (.I0(\r3_reg_n_0_[4] ),
        .I1(\r2_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_13 
       (.I0(\r7_reg_n_0_[4] ),
        .I1(\r6_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[4]_inst_i_2 
       (.I0(\RD1_OBUF[4]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[4]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[4]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[4]_inst_i_3 
       (.I0(\RD1_OBUF[4]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[4]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[4]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[4]_inst_i_4 
       (.I0(\RD1_OBUF[4]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[4]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[4]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[4]_inst_i_5 
       (.I0(\RD1_OBUF[4]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[4]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[4]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_6 
       (.I0(\r27_reg_n_0_[4] ),
        .I1(\r26_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_7 
       (.I0(\r31_reg_n_0_[4] ),
        .I1(\r30_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_8 
       (.I0(\r19_reg_n_0_[4] ),
        .I1(\r18_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[4]_inst_i_9 
       (.I0(\r23_reg_n_0_[4] ),
        .I1(\r22_reg_n_0_[4] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[4] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[4] ),
        .O(\RD1_OBUF[4]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[5]_inst 
       (.I(RD1_OBUF[5]),
        .O(RD1[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_1 
       (.I0(\RD1_OBUF[5]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[5]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[5]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[5]_inst_i_5_n_0 ),
        .O(RD1_OBUF[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_10 
       (.I0(\r11_reg_n_0_[5] ),
        .I1(\r10_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_11 
       (.I0(\r15_reg_n_0_[5] ),
        .I1(\r14_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[5]_inst_i_12 
       (.I0(\r3_reg_n_0_[5] ),
        .I1(\r2_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_13 
       (.I0(\r7_reg_n_0_[5] ),
        .I1(\r6_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[5]_inst_i_2 
       (.I0(\RD1_OBUF[5]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[5]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[5]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[5]_inst_i_3 
       (.I0(\RD1_OBUF[5]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[5]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[5]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[5]_inst_i_4 
       (.I0(\RD1_OBUF[5]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[5]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[5]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[5]_inst_i_5 
       (.I0(\RD1_OBUF[5]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[5]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[5]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_6 
       (.I0(\r27_reg_n_0_[5] ),
        .I1(\r26_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_7 
       (.I0(\r31_reg_n_0_[5] ),
        .I1(\r30_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_8 
       (.I0(\r19_reg_n_0_[5] ),
        .I1(\r18_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[5]_inst_i_9 
       (.I0(\r23_reg_n_0_[5] ),
        .I1(\r22_reg_n_0_[5] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[5] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[5] ),
        .O(\RD1_OBUF[5]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[6]_inst 
       (.I(RD1_OBUF[6]),
        .O(RD1[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_1 
       (.I0(\RD1_OBUF[6]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[6]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[6]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[6]_inst_i_5_n_0 ),
        .O(RD1_OBUF[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_10 
       (.I0(\r11_reg_n_0_[6] ),
        .I1(\r10_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_11 
       (.I0(\r15_reg_n_0_[6] ),
        .I1(\r14_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[6]_inst_i_12 
       (.I0(\r3_reg_n_0_[6] ),
        .I1(\r2_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_13 
       (.I0(\r7_reg_n_0_[6] ),
        .I1(\r6_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[6]_inst_i_2 
       (.I0(\RD1_OBUF[6]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[6]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[6]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[6]_inst_i_3 
       (.I0(\RD1_OBUF[6]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[6]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[6]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[6]_inst_i_4 
       (.I0(\RD1_OBUF[6]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[6]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[6]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[6]_inst_i_5 
       (.I0(\RD1_OBUF[6]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[6]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[6]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_6 
       (.I0(\r27_reg_n_0_[6] ),
        .I1(\r26_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_7 
       (.I0(\r31_reg_n_0_[6] ),
        .I1(\r30_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_8 
       (.I0(\r19_reg_n_0_[6] ),
        .I1(\r18_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[6]_inst_i_9 
       (.I0(\r23_reg_n_0_[6] ),
        .I1(\r22_reg_n_0_[6] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[6] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[6] ),
        .O(\RD1_OBUF[6]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[7]_inst 
       (.I(RD1_OBUF[7]),
        .O(RD1[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_1 
       (.I0(\RD1_OBUF[7]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[7]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[7]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[7]_inst_i_5_n_0 ),
        .O(RD1_OBUF[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_10 
       (.I0(\r11_reg_n_0_[7] ),
        .I1(\r10_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_11 
       (.I0(\r15_reg_n_0_[7] ),
        .I1(\r14_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[7]_inst_i_12 
       (.I0(\r3_reg_n_0_[7] ),
        .I1(\r2_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_13 
       (.I0(\r7_reg_n_0_[7] ),
        .I1(\r6_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[7]_inst_i_2 
       (.I0(\RD1_OBUF[7]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[7]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[7]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[7]_inst_i_3 
       (.I0(\RD1_OBUF[7]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[7]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[7]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[7]_inst_i_4 
       (.I0(\RD1_OBUF[7]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[7]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[7]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[7]_inst_i_5 
       (.I0(\RD1_OBUF[7]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[7]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[7]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_6 
       (.I0(\r27_reg_n_0_[7] ),
        .I1(\r26_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_7 
       (.I0(\r31_reg_n_0_[7] ),
        .I1(\r30_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_8 
       (.I0(\r19_reg_n_0_[7] ),
        .I1(\r18_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[7]_inst_i_9 
       (.I0(\r23_reg_n_0_[7] ),
        .I1(\r22_reg_n_0_[7] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[7] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[7] ),
        .O(\RD1_OBUF[7]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[8]_inst 
       (.I(RD1_OBUF[8]),
        .O(RD1[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_1 
       (.I0(\RD1_OBUF[8]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[8]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[8]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[8]_inst_i_5_n_0 ),
        .O(RD1_OBUF[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_10 
       (.I0(\r11_reg_n_0_[8] ),
        .I1(\r10_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_11 
       (.I0(\r15_reg_n_0_[8] ),
        .I1(\r14_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[8]_inst_i_12 
       (.I0(\r3_reg_n_0_[8] ),
        .I1(\r2_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_13 
       (.I0(\r7_reg_n_0_[8] ),
        .I1(\r6_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[8]_inst_i_2 
       (.I0(\RD1_OBUF[8]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[8]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[8]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[8]_inst_i_3 
       (.I0(\RD1_OBUF[8]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[8]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[8]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[8]_inst_i_4 
       (.I0(\RD1_OBUF[8]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[8]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[8]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[8]_inst_i_5 
       (.I0(\RD1_OBUF[8]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[8]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[8]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_6 
       (.I0(\r27_reg_n_0_[8] ),
        .I1(\r26_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_7 
       (.I0(\r31_reg_n_0_[8] ),
        .I1(\r30_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_8 
       (.I0(\r19_reg_n_0_[8] ),
        .I1(\r18_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[8]_inst_i_9 
       (.I0(\r23_reg_n_0_[8] ),
        .I1(\r22_reg_n_0_[8] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[8] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[8] ),
        .O(\RD1_OBUF[8]_inst_i_9_n_0 ));
  OBUF \RD1_OBUF[9]_inst 
       (.I(RD1_OBUF[9]),
        .O(RD1[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_1 
       (.I0(\RD1_OBUF[9]_inst_i_2_n_0 ),
        .I1(\RD1_OBUF[9]_inst_i_3_n_0 ),
        .I2(A1_IBUF[4]),
        .I3(\RD1_OBUF[9]_inst_i_4_n_0 ),
        .I4(A1_IBUF[3]),
        .I5(\RD1_OBUF[9]_inst_i_5_n_0 ),
        .O(RD1_OBUF[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_10 
       (.I0(\r11_reg_n_0_[9] ),
        .I1(\r10_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r9_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r8_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_11 
       (.I0(\r15_reg_n_0_[9] ),
        .I1(\r14_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r13_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r12_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD1_OBUF[9]_inst_i_12 
       (.I0(\r3_reg_n_0_[9] ),
        .I1(\r2_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(A1_IBUF[0]),
        .I4(\r1_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_13 
       (.I0(\r7_reg_n_0_[9] ),
        .I1(\r6_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r5_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r4_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_13_n_0 ));
  MUXF7 \RD1_OBUF[9]_inst_i_2 
       (.I0(\RD1_OBUF[9]_inst_i_6_n_0 ),
        .I1(\RD1_OBUF[9]_inst_i_7_n_0 ),
        .O(\RD1_OBUF[9]_inst_i_2_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[9]_inst_i_3 
       (.I0(\RD1_OBUF[9]_inst_i_8_n_0 ),
        .I1(\RD1_OBUF[9]_inst_i_9_n_0 ),
        .O(\RD1_OBUF[9]_inst_i_3_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[9]_inst_i_4 
       (.I0(\RD1_OBUF[9]_inst_i_10_n_0 ),
        .I1(\RD1_OBUF[9]_inst_i_11_n_0 ),
        .O(\RD1_OBUF[9]_inst_i_4_n_0 ),
        .S(A1_IBUF[2]));
  MUXF7 \RD1_OBUF[9]_inst_i_5 
       (.I0(\RD1_OBUF[9]_inst_i_12_n_0 ),
        .I1(\RD1_OBUF[9]_inst_i_13_n_0 ),
        .O(\RD1_OBUF[9]_inst_i_5_n_0 ),
        .S(A1_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_6 
       (.I0(\r27_reg_n_0_[9] ),
        .I1(\r26_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r25_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r24_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_7 
       (.I0(\r31_reg_n_0_[9] ),
        .I1(\r30_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r29_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r28_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_8 
       (.I0(\r19_reg_n_0_[9] ),
        .I1(\r18_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r17_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r16_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD1_OBUF[9]_inst_i_9 
       (.I0(\r23_reg_n_0_[9] ),
        .I1(\r22_reg_n_0_[9] ),
        .I2(A1_IBUF[1]),
        .I3(\r21_reg_n_0_[9] ),
        .I4(A1_IBUF[0]),
        .I5(\r20_reg_n_0_[9] ),
        .O(\RD1_OBUF[9]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[0]_inst 
       (.I(RD2_OBUF[0]),
        .O(RD2[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_1 
       (.I0(\RD2_OBUF[0]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[0]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[0]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[0]_inst_i_5_n_0 ),
        .O(RD2_OBUF[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_10 
       (.I0(\r11_reg_n_0_[0] ),
        .I1(\r10_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_11 
       (.I0(\r15_reg_n_0_[0] ),
        .I1(\r14_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[0]_inst_i_12 
       (.I0(\r3_reg_n_0_[0] ),
        .I1(\r2_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_13 
       (.I0(\r7_reg_n_0_[0] ),
        .I1(\r6_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[0]_inst_i_2 
       (.I0(\RD2_OBUF[0]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[0]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[0]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[0]_inst_i_3 
       (.I0(\RD2_OBUF[0]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[0]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[0]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[0]_inst_i_4 
       (.I0(\RD2_OBUF[0]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[0]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[0]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[0]_inst_i_5 
       (.I0(\RD2_OBUF[0]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[0]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[0]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_6 
       (.I0(\r27_reg_n_0_[0] ),
        .I1(\r26_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_7 
       (.I0(\r31_reg_n_0_[0] ),
        .I1(\r30_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_8 
       (.I0(\r19_reg_n_0_[0] ),
        .I1(\r18_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[0]_inst_i_9 
       (.I0(\r23_reg_n_0_[0] ),
        .I1(\r22_reg_n_0_[0] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[0] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[0] ),
        .O(\RD2_OBUF[0]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[10]_inst 
       (.I(RD2_OBUF[10]),
        .O(RD2[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_1 
       (.I0(\RD2_OBUF[10]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[10]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[10]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[10]_inst_i_5_n_0 ),
        .O(RD2_OBUF[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_10 
       (.I0(\r11_reg_n_0_[10] ),
        .I1(\r10_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_11 
       (.I0(\r15_reg_n_0_[10] ),
        .I1(\r14_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[10]_inst_i_12 
       (.I0(\r3_reg_n_0_[10] ),
        .I1(\r2_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_13 
       (.I0(\r7_reg_n_0_[10] ),
        .I1(\r6_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[10]_inst_i_2 
       (.I0(\RD2_OBUF[10]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[10]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[10]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[10]_inst_i_3 
       (.I0(\RD2_OBUF[10]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[10]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[10]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[10]_inst_i_4 
       (.I0(\RD2_OBUF[10]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[10]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[10]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[10]_inst_i_5 
       (.I0(\RD2_OBUF[10]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[10]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[10]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_6 
       (.I0(\r27_reg_n_0_[10] ),
        .I1(\r26_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_7 
       (.I0(\r31_reg_n_0_[10] ),
        .I1(\r30_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_8 
       (.I0(\r19_reg_n_0_[10] ),
        .I1(\r18_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[10]_inst_i_9 
       (.I0(\r23_reg_n_0_[10] ),
        .I1(\r22_reg_n_0_[10] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[10] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[10] ),
        .O(\RD2_OBUF[10]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[11]_inst 
       (.I(RD2_OBUF[11]),
        .O(RD2[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_1 
       (.I0(\RD2_OBUF[11]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[11]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[11]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[11]_inst_i_5_n_0 ),
        .O(RD2_OBUF[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_10 
       (.I0(\r11_reg_n_0_[11] ),
        .I1(\r10_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_11 
       (.I0(\r15_reg_n_0_[11] ),
        .I1(\r14_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[11]_inst_i_12 
       (.I0(\r3_reg_n_0_[11] ),
        .I1(\r2_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_13 
       (.I0(\r7_reg_n_0_[11] ),
        .I1(\r6_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[11]_inst_i_2 
       (.I0(\RD2_OBUF[11]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[11]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[11]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[11]_inst_i_3 
       (.I0(\RD2_OBUF[11]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[11]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[11]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[11]_inst_i_4 
       (.I0(\RD2_OBUF[11]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[11]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[11]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[11]_inst_i_5 
       (.I0(\RD2_OBUF[11]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[11]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[11]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_6 
       (.I0(\r27_reg_n_0_[11] ),
        .I1(\r26_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_7 
       (.I0(\r31_reg_n_0_[11] ),
        .I1(\r30_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_8 
       (.I0(\r19_reg_n_0_[11] ),
        .I1(\r18_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[11]_inst_i_9 
       (.I0(\r23_reg_n_0_[11] ),
        .I1(\r22_reg_n_0_[11] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[11] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[11] ),
        .O(\RD2_OBUF[11]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[12]_inst 
       (.I(RD2_OBUF[12]),
        .O(RD2[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_1 
       (.I0(\RD2_OBUF[12]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[12]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[12]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[12]_inst_i_5_n_0 ),
        .O(RD2_OBUF[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_10 
       (.I0(\r11_reg_n_0_[12] ),
        .I1(\r10_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_11 
       (.I0(\r15_reg_n_0_[12] ),
        .I1(\r14_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[12]_inst_i_12 
       (.I0(\r3_reg_n_0_[12] ),
        .I1(\r2_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_13 
       (.I0(\r7_reg_n_0_[12] ),
        .I1(\r6_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[12]_inst_i_2 
       (.I0(\RD2_OBUF[12]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[12]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[12]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[12]_inst_i_3 
       (.I0(\RD2_OBUF[12]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[12]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[12]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[12]_inst_i_4 
       (.I0(\RD2_OBUF[12]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[12]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[12]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[12]_inst_i_5 
       (.I0(\RD2_OBUF[12]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[12]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[12]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_6 
       (.I0(\r27_reg_n_0_[12] ),
        .I1(\r26_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_7 
       (.I0(\r31_reg_n_0_[12] ),
        .I1(\r30_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_8 
       (.I0(\r19_reg_n_0_[12] ),
        .I1(\r18_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[12]_inst_i_9 
       (.I0(\r23_reg_n_0_[12] ),
        .I1(\r22_reg_n_0_[12] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[12] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[12] ),
        .O(\RD2_OBUF[12]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[13]_inst 
       (.I(RD2_OBUF[13]),
        .O(RD2[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_1 
       (.I0(\RD2_OBUF[13]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[13]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[13]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[13]_inst_i_5_n_0 ),
        .O(RD2_OBUF[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_10 
       (.I0(\r11_reg_n_0_[13] ),
        .I1(\r10_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_11 
       (.I0(\r15_reg_n_0_[13] ),
        .I1(\r14_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[13]_inst_i_12 
       (.I0(\r3_reg_n_0_[13] ),
        .I1(\r2_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_13 
       (.I0(\r7_reg_n_0_[13] ),
        .I1(\r6_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[13]_inst_i_2 
       (.I0(\RD2_OBUF[13]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[13]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[13]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[13]_inst_i_3 
       (.I0(\RD2_OBUF[13]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[13]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[13]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[13]_inst_i_4 
       (.I0(\RD2_OBUF[13]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[13]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[13]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[13]_inst_i_5 
       (.I0(\RD2_OBUF[13]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[13]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[13]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_6 
       (.I0(\r27_reg_n_0_[13] ),
        .I1(\r26_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_7 
       (.I0(\r31_reg_n_0_[13] ),
        .I1(\r30_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_8 
       (.I0(\r19_reg_n_0_[13] ),
        .I1(\r18_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[13]_inst_i_9 
       (.I0(\r23_reg_n_0_[13] ),
        .I1(\r22_reg_n_0_[13] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[13] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[13] ),
        .O(\RD2_OBUF[13]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[14]_inst 
       (.I(RD2_OBUF[14]),
        .O(RD2[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_1 
       (.I0(\RD2_OBUF[14]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[14]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[14]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[14]_inst_i_5_n_0 ),
        .O(RD2_OBUF[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_10 
       (.I0(\r11_reg_n_0_[14] ),
        .I1(\r10_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_11 
       (.I0(\r15_reg_n_0_[14] ),
        .I1(\r14_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[14]_inst_i_12 
       (.I0(\r3_reg_n_0_[14] ),
        .I1(\r2_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_13 
       (.I0(\r7_reg_n_0_[14] ),
        .I1(\r6_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[14]_inst_i_2 
       (.I0(\RD2_OBUF[14]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[14]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[14]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[14]_inst_i_3 
       (.I0(\RD2_OBUF[14]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[14]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[14]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[14]_inst_i_4 
       (.I0(\RD2_OBUF[14]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[14]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[14]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[14]_inst_i_5 
       (.I0(\RD2_OBUF[14]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[14]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[14]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_6 
       (.I0(\r27_reg_n_0_[14] ),
        .I1(\r26_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_7 
       (.I0(\r31_reg_n_0_[14] ),
        .I1(\r30_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_8 
       (.I0(\r19_reg_n_0_[14] ),
        .I1(\r18_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[14]_inst_i_9 
       (.I0(\r23_reg_n_0_[14] ),
        .I1(\r22_reg_n_0_[14] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[14] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[14] ),
        .O(\RD2_OBUF[14]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[15]_inst 
       (.I(RD2_OBUF[15]),
        .O(RD2[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_1 
       (.I0(\RD2_OBUF[15]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[15]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[15]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[15]_inst_i_5_n_0 ),
        .O(RD2_OBUF[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_10 
       (.I0(\r11_reg_n_0_[15] ),
        .I1(\r10_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_11 
       (.I0(\r15_reg_n_0_[15] ),
        .I1(\r14_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[15]_inst_i_12 
       (.I0(\r3_reg_n_0_[15] ),
        .I1(\r2_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_13 
       (.I0(\r7_reg_n_0_[15] ),
        .I1(\r6_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[15]_inst_i_2 
       (.I0(\RD2_OBUF[15]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[15]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[15]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[15]_inst_i_3 
       (.I0(\RD2_OBUF[15]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[15]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[15]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[15]_inst_i_4 
       (.I0(\RD2_OBUF[15]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[15]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[15]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[15]_inst_i_5 
       (.I0(\RD2_OBUF[15]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[15]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[15]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_6 
       (.I0(\r27_reg_n_0_[15] ),
        .I1(\r26_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_7 
       (.I0(\r31_reg_n_0_[15] ),
        .I1(\r30_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_8 
       (.I0(\r19_reg_n_0_[15] ),
        .I1(\r18_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[15]_inst_i_9 
       (.I0(\r23_reg_n_0_[15] ),
        .I1(\r22_reg_n_0_[15] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[15] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[15] ),
        .O(\RD2_OBUF[15]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[16]_inst 
       (.I(RD2_OBUF[16]),
        .O(RD2[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_1 
       (.I0(\RD2_OBUF[16]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[16]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[16]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[16]_inst_i_5_n_0 ),
        .O(RD2_OBUF[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_10 
       (.I0(\r11_reg_n_0_[16] ),
        .I1(\r10_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_11 
       (.I0(\r15_reg_n_0_[16] ),
        .I1(\r14_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[16]_inst_i_12 
       (.I0(\r3_reg_n_0_[16] ),
        .I1(\r2_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_13 
       (.I0(\r7_reg_n_0_[16] ),
        .I1(\r6_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[16]_inst_i_2 
       (.I0(\RD2_OBUF[16]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[16]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[16]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[16]_inst_i_3 
       (.I0(\RD2_OBUF[16]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[16]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[16]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[16]_inst_i_4 
       (.I0(\RD2_OBUF[16]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[16]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[16]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[16]_inst_i_5 
       (.I0(\RD2_OBUF[16]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[16]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[16]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_6 
       (.I0(\r27_reg_n_0_[16] ),
        .I1(\r26_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_7 
       (.I0(\r31_reg_n_0_[16] ),
        .I1(\r30_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_8 
       (.I0(\r19_reg_n_0_[16] ),
        .I1(\r18_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[16]_inst_i_9 
       (.I0(\r23_reg_n_0_[16] ),
        .I1(\r22_reg_n_0_[16] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[16] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[16] ),
        .O(\RD2_OBUF[16]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[17]_inst 
       (.I(RD2_OBUF[17]),
        .O(RD2[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_1 
       (.I0(\RD2_OBUF[17]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[17]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[17]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[17]_inst_i_5_n_0 ),
        .O(RD2_OBUF[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_10 
       (.I0(\r11_reg_n_0_[17] ),
        .I1(\r10_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_11 
       (.I0(\r15_reg_n_0_[17] ),
        .I1(\r14_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[17]_inst_i_12 
       (.I0(\r3_reg_n_0_[17] ),
        .I1(\r2_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_13 
       (.I0(\r7_reg_n_0_[17] ),
        .I1(\r6_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[17]_inst_i_2 
       (.I0(\RD2_OBUF[17]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[17]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[17]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[17]_inst_i_3 
       (.I0(\RD2_OBUF[17]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[17]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[17]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[17]_inst_i_4 
       (.I0(\RD2_OBUF[17]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[17]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[17]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[17]_inst_i_5 
       (.I0(\RD2_OBUF[17]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[17]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[17]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_6 
       (.I0(\r27_reg_n_0_[17] ),
        .I1(\r26_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_7 
       (.I0(\r31_reg_n_0_[17] ),
        .I1(\r30_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_8 
       (.I0(\r19_reg_n_0_[17] ),
        .I1(\r18_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[17]_inst_i_9 
       (.I0(\r23_reg_n_0_[17] ),
        .I1(\r22_reg_n_0_[17] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[17] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[17] ),
        .O(\RD2_OBUF[17]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[18]_inst 
       (.I(RD2_OBUF[18]),
        .O(RD2[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_1 
       (.I0(\RD2_OBUF[18]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[18]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[18]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[18]_inst_i_5_n_0 ),
        .O(RD2_OBUF[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_10 
       (.I0(\r11_reg_n_0_[18] ),
        .I1(\r10_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_11 
       (.I0(\r15_reg_n_0_[18] ),
        .I1(\r14_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[18]_inst_i_12 
       (.I0(\r3_reg_n_0_[18] ),
        .I1(\r2_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_13 
       (.I0(\r7_reg_n_0_[18] ),
        .I1(\r6_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[18]_inst_i_2 
       (.I0(\RD2_OBUF[18]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[18]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[18]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[18]_inst_i_3 
       (.I0(\RD2_OBUF[18]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[18]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[18]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[18]_inst_i_4 
       (.I0(\RD2_OBUF[18]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[18]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[18]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[18]_inst_i_5 
       (.I0(\RD2_OBUF[18]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[18]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[18]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_6 
       (.I0(\r27_reg_n_0_[18] ),
        .I1(\r26_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_7 
       (.I0(\r31_reg_n_0_[18] ),
        .I1(\r30_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_8 
       (.I0(\r19_reg_n_0_[18] ),
        .I1(\r18_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[18]_inst_i_9 
       (.I0(\r23_reg_n_0_[18] ),
        .I1(\r22_reg_n_0_[18] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[18] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[18] ),
        .O(\RD2_OBUF[18]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[19]_inst 
       (.I(RD2_OBUF[19]),
        .O(RD2[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_1 
       (.I0(\RD2_OBUF[19]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[19]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[19]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[19]_inst_i_5_n_0 ),
        .O(RD2_OBUF[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_10 
       (.I0(\r11_reg_n_0_[19] ),
        .I1(\r10_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_11 
       (.I0(\r15_reg_n_0_[19] ),
        .I1(\r14_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[19]_inst_i_12 
       (.I0(\r3_reg_n_0_[19] ),
        .I1(\r2_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_13 
       (.I0(\r7_reg_n_0_[19] ),
        .I1(\r6_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[19]_inst_i_2 
       (.I0(\RD2_OBUF[19]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[19]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[19]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[19]_inst_i_3 
       (.I0(\RD2_OBUF[19]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[19]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[19]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[19]_inst_i_4 
       (.I0(\RD2_OBUF[19]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[19]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[19]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[19]_inst_i_5 
       (.I0(\RD2_OBUF[19]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[19]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[19]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_6 
       (.I0(\r27_reg_n_0_[19] ),
        .I1(\r26_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_7 
       (.I0(\r31_reg_n_0_[19] ),
        .I1(\r30_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_8 
       (.I0(\r19_reg_n_0_[19] ),
        .I1(\r18_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[19]_inst_i_9 
       (.I0(\r23_reg_n_0_[19] ),
        .I1(\r22_reg_n_0_[19] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[19] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[19] ),
        .O(\RD2_OBUF[19]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[1]_inst 
       (.I(RD2_OBUF[1]),
        .O(RD2[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_1 
       (.I0(\RD2_OBUF[1]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[1]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[1]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[1]_inst_i_5_n_0 ),
        .O(RD2_OBUF[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_10 
       (.I0(\r11_reg_n_0_[1] ),
        .I1(\r10_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_11 
       (.I0(\r15_reg_n_0_[1] ),
        .I1(\r14_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[1]_inst_i_12 
       (.I0(\r3_reg_n_0_[1] ),
        .I1(\r2_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_13 
       (.I0(\r7_reg_n_0_[1] ),
        .I1(\r6_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[1]_inst_i_2 
       (.I0(\RD2_OBUF[1]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[1]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[1]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[1]_inst_i_3 
       (.I0(\RD2_OBUF[1]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[1]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[1]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[1]_inst_i_4 
       (.I0(\RD2_OBUF[1]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[1]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[1]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[1]_inst_i_5 
       (.I0(\RD2_OBUF[1]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[1]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[1]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_6 
       (.I0(\r27_reg_n_0_[1] ),
        .I1(\r26_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_7 
       (.I0(\r31_reg_n_0_[1] ),
        .I1(\r30_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_8 
       (.I0(\r19_reg_n_0_[1] ),
        .I1(\r18_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[1]_inst_i_9 
       (.I0(\r23_reg_n_0_[1] ),
        .I1(\r22_reg_n_0_[1] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[1] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[1] ),
        .O(\RD2_OBUF[1]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[20]_inst 
       (.I(RD2_OBUF[20]),
        .O(RD2[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_1 
       (.I0(\RD2_OBUF[20]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[20]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[20]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[20]_inst_i_5_n_0 ),
        .O(RD2_OBUF[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_10 
       (.I0(\r11_reg_n_0_[20] ),
        .I1(\r10_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_11 
       (.I0(\r15_reg_n_0_[20] ),
        .I1(\r14_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[20]_inst_i_12 
       (.I0(\r3_reg_n_0_[20] ),
        .I1(\r2_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_13 
       (.I0(\r7_reg_n_0_[20] ),
        .I1(\r6_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[20]_inst_i_2 
       (.I0(\RD2_OBUF[20]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[20]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[20]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[20]_inst_i_3 
       (.I0(\RD2_OBUF[20]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[20]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[20]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[20]_inst_i_4 
       (.I0(\RD2_OBUF[20]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[20]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[20]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[20]_inst_i_5 
       (.I0(\RD2_OBUF[20]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[20]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[20]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_6 
       (.I0(\r27_reg_n_0_[20] ),
        .I1(\r26_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_7 
       (.I0(\r31_reg_n_0_[20] ),
        .I1(\r30_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_8 
       (.I0(\r19_reg_n_0_[20] ),
        .I1(\r18_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[20]_inst_i_9 
       (.I0(\r23_reg_n_0_[20] ),
        .I1(\r22_reg_n_0_[20] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[20] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[20] ),
        .O(\RD2_OBUF[20]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[21]_inst 
       (.I(RD2_OBUF[21]),
        .O(RD2[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_1 
       (.I0(\RD2_OBUF[21]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[21]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[21]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[21]_inst_i_5_n_0 ),
        .O(RD2_OBUF[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_10 
       (.I0(\r11_reg_n_0_[21] ),
        .I1(\r10_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_11 
       (.I0(\r15_reg_n_0_[21] ),
        .I1(\r14_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[21]_inst_i_12 
       (.I0(\r3_reg_n_0_[21] ),
        .I1(\r2_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_13 
       (.I0(\r7_reg_n_0_[21] ),
        .I1(\r6_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[21]_inst_i_2 
       (.I0(\RD2_OBUF[21]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[21]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[21]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[21]_inst_i_3 
       (.I0(\RD2_OBUF[21]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[21]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[21]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[21]_inst_i_4 
       (.I0(\RD2_OBUF[21]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[21]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[21]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[21]_inst_i_5 
       (.I0(\RD2_OBUF[21]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[21]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[21]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_6 
       (.I0(\r27_reg_n_0_[21] ),
        .I1(\r26_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_7 
       (.I0(\r31_reg_n_0_[21] ),
        .I1(\r30_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_8 
       (.I0(\r19_reg_n_0_[21] ),
        .I1(\r18_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[21]_inst_i_9 
       (.I0(\r23_reg_n_0_[21] ),
        .I1(\r22_reg_n_0_[21] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[21] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[21] ),
        .O(\RD2_OBUF[21]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[22]_inst 
       (.I(RD2_OBUF[22]),
        .O(RD2[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_1 
       (.I0(\RD2_OBUF[22]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[22]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[22]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[22]_inst_i_5_n_0 ),
        .O(RD2_OBUF[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_10 
       (.I0(\r11_reg_n_0_[22] ),
        .I1(\r10_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_11 
       (.I0(\r15_reg_n_0_[22] ),
        .I1(\r14_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[22]_inst_i_12 
       (.I0(\r3_reg_n_0_[22] ),
        .I1(\r2_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_13 
       (.I0(\r7_reg_n_0_[22] ),
        .I1(\r6_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[22]_inst_i_2 
       (.I0(\RD2_OBUF[22]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[22]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[22]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[22]_inst_i_3 
       (.I0(\RD2_OBUF[22]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[22]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[22]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[22]_inst_i_4 
       (.I0(\RD2_OBUF[22]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[22]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[22]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[22]_inst_i_5 
       (.I0(\RD2_OBUF[22]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[22]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[22]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_6 
       (.I0(\r27_reg_n_0_[22] ),
        .I1(\r26_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_7 
       (.I0(\r31_reg_n_0_[22] ),
        .I1(\r30_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_8 
       (.I0(\r19_reg_n_0_[22] ),
        .I1(\r18_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[22]_inst_i_9 
       (.I0(\r23_reg_n_0_[22] ),
        .I1(\r22_reg_n_0_[22] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[22] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[22] ),
        .O(\RD2_OBUF[22]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[23]_inst 
       (.I(RD2_OBUF[23]),
        .O(RD2[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_1 
       (.I0(\RD2_OBUF[23]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[23]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[23]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[23]_inst_i_5_n_0 ),
        .O(RD2_OBUF[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_10 
       (.I0(\r11_reg_n_0_[23] ),
        .I1(\r10_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_11 
       (.I0(\r15_reg_n_0_[23] ),
        .I1(\r14_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[23]_inst_i_12 
       (.I0(\r3_reg_n_0_[23] ),
        .I1(\r2_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_13 
       (.I0(\r7_reg_n_0_[23] ),
        .I1(\r6_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[23]_inst_i_2 
       (.I0(\RD2_OBUF[23]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[23]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[23]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[23]_inst_i_3 
       (.I0(\RD2_OBUF[23]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[23]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[23]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[23]_inst_i_4 
       (.I0(\RD2_OBUF[23]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[23]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[23]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[23]_inst_i_5 
       (.I0(\RD2_OBUF[23]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[23]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[23]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_6 
       (.I0(\r27_reg_n_0_[23] ),
        .I1(\r26_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_7 
       (.I0(\r31_reg_n_0_[23] ),
        .I1(\r30_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_8 
       (.I0(\r19_reg_n_0_[23] ),
        .I1(\r18_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[23]_inst_i_9 
       (.I0(\r23_reg_n_0_[23] ),
        .I1(\r22_reg_n_0_[23] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[23] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[23] ),
        .O(\RD2_OBUF[23]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[24]_inst 
       (.I(RD2_OBUF[24]),
        .O(RD2[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_1 
       (.I0(\RD2_OBUF[24]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[24]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[24]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[24]_inst_i_5_n_0 ),
        .O(RD2_OBUF[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_10 
       (.I0(\r11_reg_n_0_[24] ),
        .I1(\r10_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_11 
       (.I0(\r15_reg_n_0_[24] ),
        .I1(\r14_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[24]_inst_i_12 
       (.I0(\r3_reg_n_0_[24] ),
        .I1(\r2_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_13 
       (.I0(\r7_reg_n_0_[24] ),
        .I1(\r6_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[24]_inst_i_2 
       (.I0(\RD2_OBUF[24]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[24]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[24]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[24]_inst_i_3 
       (.I0(\RD2_OBUF[24]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[24]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[24]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[24]_inst_i_4 
       (.I0(\RD2_OBUF[24]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[24]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[24]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[24]_inst_i_5 
       (.I0(\RD2_OBUF[24]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[24]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[24]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_6 
       (.I0(\r27_reg_n_0_[24] ),
        .I1(\r26_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_7 
       (.I0(\r31_reg_n_0_[24] ),
        .I1(\r30_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_8 
       (.I0(\r19_reg_n_0_[24] ),
        .I1(\r18_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[24]_inst_i_9 
       (.I0(\r23_reg_n_0_[24] ),
        .I1(\r22_reg_n_0_[24] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[24] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[24] ),
        .O(\RD2_OBUF[24]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[25]_inst 
       (.I(RD2_OBUF[25]),
        .O(RD2[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_1 
       (.I0(\RD2_OBUF[25]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[25]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[25]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[25]_inst_i_5_n_0 ),
        .O(RD2_OBUF[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_10 
       (.I0(\r11_reg_n_0_[25] ),
        .I1(\r10_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_11 
       (.I0(\r15_reg_n_0_[25] ),
        .I1(\r14_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[25]_inst_i_12 
       (.I0(\r3_reg_n_0_[25] ),
        .I1(\r2_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_13 
       (.I0(\r7_reg_n_0_[25] ),
        .I1(\r6_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[25]_inst_i_2 
       (.I0(\RD2_OBUF[25]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[25]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[25]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[25]_inst_i_3 
       (.I0(\RD2_OBUF[25]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[25]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[25]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[25]_inst_i_4 
       (.I0(\RD2_OBUF[25]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[25]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[25]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[25]_inst_i_5 
       (.I0(\RD2_OBUF[25]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[25]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[25]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_6 
       (.I0(\r27_reg_n_0_[25] ),
        .I1(\r26_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_7 
       (.I0(\r31_reg_n_0_[25] ),
        .I1(\r30_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_8 
       (.I0(\r19_reg_n_0_[25] ),
        .I1(\r18_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[25]_inst_i_9 
       (.I0(\r23_reg_n_0_[25] ),
        .I1(\r22_reg_n_0_[25] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[25] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[25] ),
        .O(\RD2_OBUF[25]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[26]_inst 
       (.I(RD2_OBUF[26]),
        .O(RD2[26]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_1 
       (.I0(\RD2_OBUF[26]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[26]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[26]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[26]_inst_i_5_n_0 ),
        .O(RD2_OBUF[26]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_10 
       (.I0(\r11_reg_n_0_[26] ),
        .I1(\r10_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_11 
       (.I0(\r15_reg_n_0_[26] ),
        .I1(\r14_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[26]_inst_i_12 
       (.I0(\r3_reg_n_0_[26] ),
        .I1(\r2_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_13 
       (.I0(\r7_reg_n_0_[26] ),
        .I1(\r6_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[26]_inst_i_2 
       (.I0(\RD2_OBUF[26]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[26]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[26]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[26]_inst_i_3 
       (.I0(\RD2_OBUF[26]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[26]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[26]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[26]_inst_i_4 
       (.I0(\RD2_OBUF[26]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[26]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[26]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[26]_inst_i_5 
       (.I0(\RD2_OBUF[26]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[26]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[26]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_6 
       (.I0(\r27_reg_n_0_[26] ),
        .I1(\r26_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_7 
       (.I0(\r31_reg_n_0_[26] ),
        .I1(\r30_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_8 
       (.I0(\r19_reg_n_0_[26] ),
        .I1(\r18_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[26]_inst_i_9 
       (.I0(\r23_reg_n_0_[26] ),
        .I1(\r22_reg_n_0_[26] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[26] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[26] ),
        .O(\RD2_OBUF[26]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[27]_inst 
       (.I(RD2_OBUF[27]),
        .O(RD2[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_1 
       (.I0(\RD2_OBUF[27]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[27]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[27]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[27]_inst_i_5_n_0 ),
        .O(RD2_OBUF[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_10 
       (.I0(\r11_reg_n_0_[27] ),
        .I1(\r10_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_11 
       (.I0(\r15_reg_n_0_[27] ),
        .I1(\r14_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[27]_inst_i_12 
       (.I0(\r3_reg_n_0_[27] ),
        .I1(\r2_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_13 
       (.I0(\r7_reg_n_0_[27] ),
        .I1(\r6_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[27]_inst_i_2 
       (.I0(\RD2_OBUF[27]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[27]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[27]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[27]_inst_i_3 
       (.I0(\RD2_OBUF[27]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[27]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[27]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[27]_inst_i_4 
       (.I0(\RD2_OBUF[27]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[27]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[27]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[27]_inst_i_5 
       (.I0(\RD2_OBUF[27]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[27]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[27]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_6 
       (.I0(\r27_reg_n_0_[27] ),
        .I1(\r26_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_7 
       (.I0(\r31_reg_n_0_[27] ),
        .I1(\r30_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_8 
       (.I0(\r19_reg_n_0_[27] ),
        .I1(\r18_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[27]_inst_i_9 
       (.I0(\r23_reg_n_0_[27] ),
        .I1(\r22_reg_n_0_[27] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[27] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[27] ),
        .O(\RD2_OBUF[27]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[28]_inst 
       (.I(RD2_OBUF[28]),
        .O(RD2[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_1 
       (.I0(\RD2_OBUF[28]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[28]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[28]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[28]_inst_i_5_n_0 ),
        .O(RD2_OBUF[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_10 
       (.I0(\r11_reg_n_0_[28] ),
        .I1(\r10_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_11 
       (.I0(\r15_reg_n_0_[28] ),
        .I1(\r14_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[28]_inst_i_12 
       (.I0(\r3_reg_n_0_[28] ),
        .I1(\r2_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_13 
       (.I0(\r7_reg_n_0_[28] ),
        .I1(\r6_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[28]_inst_i_2 
       (.I0(\RD2_OBUF[28]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[28]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[28]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[28]_inst_i_3 
       (.I0(\RD2_OBUF[28]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[28]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[28]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[28]_inst_i_4 
       (.I0(\RD2_OBUF[28]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[28]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[28]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[28]_inst_i_5 
       (.I0(\RD2_OBUF[28]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[28]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[28]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_6 
       (.I0(\r27_reg_n_0_[28] ),
        .I1(\r26_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_7 
       (.I0(\r31_reg_n_0_[28] ),
        .I1(\r30_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_8 
       (.I0(\r19_reg_n_0_[28] ),
        .I1(\r18_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[28]_inst_i_9 
       (.I0(\r23_reg_n_0_[28] ),
        .I1(\r22_reg_n_0_[28] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[28] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[28] ),
        .O(\RD2_OBUF[28]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[29]_inst 
       (.I(RD2_OBUF[29]),
        .O(RD2[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_1 
       (.I0(\RD2_OBUF[29]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[29]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[29]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[29]_inst_i_5_n_0 ),
        .O(RD2_OBUF[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_10 
       (.I0(\r11_reg_n_0_[29] ),
        .I1(\r10_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_11 
       (.I0(\r15_reg_n_0_[29] ),
        .I1(\r14_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[29]_inst_i_12 
       (.I0(\r3_reg_n_0_[29] ),
        .I1(\r2_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_13 
       (.I0(\r7_reg_n_0_[29] ),
        .I1(\r6_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[29]_inst_i_2 
       (.I0(\RD2_OBUF[29]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[29]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[29]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[29]_inst_i_3 
       (.I0(\RD2_OBUF[29]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[29]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[29]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[29]_inst_i_4 
       (.I0(\RD2_OBUF[29]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[29]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[29]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[29]_inst_i_5 
       (.I0(\RD2_OBUF[29]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[29]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[29]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_6 
       (.I0(\r27_reg_n_0_[29] ),
        .I1(\r26_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_7 
       (.I0(\r31_reg_n_0_[29] ),
        .I1(\r30_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_8 
       (.I0(\r19_reg_n_0_[29] ),
        .I1(\r18_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[29]_inst_i_9 
       (.I0(\r23_reg_n_0_[29] ),
        .I1(\r22_reg_n_0_[29] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[29] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[29] ),
        .O(\RD2_OBUF[29]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[2]_inst 
       (.I(RD2_OBUF[2]),
        .O(RD2[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_1 
       (.I0(\RD2_OBUF[2]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[2]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[2]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[2]_inst_i_5_n_0 ),
        .O(RD2_OBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_10 
       (.I0(\r11_reg_n_0_[2] ),
        .I1(\r10_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_11 
       (.I0(\r15_reg_n_0_[2] ),
        .I1(\r14_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[2]_inst_i_12 
       (.I0(\r3_reg_n_0_[2] ),
        .I1(\r2_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_13 
       (.I0(\r7_reg_n_0_[2] ),
        .I1(\r6_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[2]_inst_i_2 
       (.I0(\RD2_OBUF[2]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[2]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[2]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[2]_inst_i_3 
       (.I0(\RD2_OBUF[2]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[2]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[2]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[2]_inst_i_4 
       (.I0(\RD2_OBUF[2]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[2]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[2]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[2]_inst_i_5 
       (.I0(\RD2_OBUF[2]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[2]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[2]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_6 
       (.I0(\r27_reg_n_0_[2] ),
        .I1(\r26_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_7 
       (.I0(\r31_reg_n_0_[2] ),
        .I1(\r30_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_8 
       (.I0(\r19_reg_n_0_[2] ),
        .I1(\r18_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[2]_inst_i_9 
       (.I0(\r23_reg_n_0_[2] ),
        .I1(\r22_reg_n_0_[2] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[2] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[2] ),
        .O(\RD2_OBUF[2]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[30]_inst 
       (.I(RD2_OBUF[30]),
        .O(RD2[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_1 
       (.I0(\RD2_OBUF[30]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[30]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[30]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[30]_inst_i_5_n_0 ),
        .O(RD2_OBUF[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_10 
       (.I0(\r11_reg_n_0_[30] ),
        .I1(\r10_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_11 
       (.I0(\r15_reg_n_0_[30] ),
        .I1(\r14_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[30]_inst_i_12 
       (.I0(\r3_reg_n_0_[30] ),
        .I1(\r2_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_13 
       (.I0(\r7_reg_n_0_[30] ),
        .I1(\r6_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[30]_inst_i_2 
       (.I0(\RD2_OBUF[30]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[30]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[30]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[30]_inst_i_3 
       (.I0(\RD2_OBUF[30]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[30]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[30]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[30]_inst_i_4 
       (.I0(\RD2_OBUF[30]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[30]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[30]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[30]_inst_i_5 
       (.I0(\RD2_OBUF[30]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[30]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[30]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_6 
       (.I0(\r27_reg_n_0_[30] ),
        .I1(\r26_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_7 
       (.I0(\r31_reg_n_0_[30] ),
        .I1(\r30_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_8 
       (.I0(\r19_reg_n_0_[30] ),
        .I1(\r18_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[30]_inst_i_9 
       (.I0(\r23_reg_n_0_[30] ),
        .I1(\r22_reg_n_0_[30] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[30] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[30] ),
        .O(\RD2_OBUF[30]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[31]_inst 
       (.I(RD2_OBUF[31]),
        .O(RD2[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_1 
       (.I0(\RD2_OBUF[31]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[31]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[31]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[31]_inst_i_5_n_0 ),
        .O(RD2_OBUF[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_10 
       (.I0(\r11_reg_n_0_[31] ),
        .I1(\r10_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_11 
       (.I0(\r15_reg_n_0_[31] ),
        .I1(\r14_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[31]_inst_i_12 
       (.I0(\r3_reg_n_0_[31] ),
        .I1(\r2_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_13 
       (.I0(\r7_reg_n_0_[31] ),
        .I1(\r6_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[31]_inst_i_2 
       (.I0(\RD2_OBUF[31]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[31]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[31]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[31]_inst_i_3 
       (.I0(\RD2_OBUF[31]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[31]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[31]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[31]_inst_i_4 
       (.I0(\RD2_OBUF[31]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[31]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[31]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[31]_inst_i_5 
       (.I0(\RD2_OBUF[31]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[31]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[31]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_6 
       (.I0(\r27_reg_n_0_[31] ),
        .I1(\r26_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_7 
       (.I0(\r31_reg_n_0_[31] ),
        .I1(\r30_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_8 
       (.I0(\r19_reg_n_0_[31] ),
        .I1(\r18_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[31]_inst_i_9 
       (.I0(\r23_reg_n_0_[31] ),
        .I1(\r22_reg_n_0_[31] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[31] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[31] ),
        .O(\RD2_OBUF[31]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[3]_inst 
       (.I(RD2_OBUF[3]),
        .O(RD2[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_1 
       (.I0(\RD2_OBUF[3]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[3]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[3]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[3]_inst_i_5_n_0 ),
        .O(RD2_OBUF[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_10 
       (.I0(\r11_reg_n_0_[3] ),
        .I1(\r10_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_11 
       (.I0(\r15_reg_n_0_[3] ),
        .I1(\r14_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[3]_inst_i_12 
       (.I0(\r3_reg_n_0_[3] ),
        .I1(\r2_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_13 
       (.I0(\r7_reg_n_0_[3] ),
        .I1(\r6_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[3]_inst_i_2 
       (.I0(\RD2_OBUF[3]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[3]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[3]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[3]_inst_i_3 
       (.I0(\RD2_OBUF[3]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[3]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[3]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[3]_inst_i_4 
       (.I0(\RD2_OBUF[3]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[3]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[3]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[3]_inst_i_5 
       (.I0(\RD2_OBUF[3]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[3]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[3]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_6 
       (.I0(\r27_reg_n_0_[3] ),
        .I1(\r26_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_7 
       (.I0(\r31_reg_n_0_[3] ),
        .I1(\r30_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_8 
       (.I0(\r19_reg_n_0_[3] ),
        .I1(\r18_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[3]_inst_i_9 
       (.I0(\r23_reg_n_0_[3] ),
        .I1(\r22_reg_n_0_[3] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[3] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[3] ),
        .O(\RD2_OBUF[3]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[4]_inst 
       (.I(RD2_OBUF[4]),
        .O(RD2[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_1 
       (.I0(\RD2_OBUF[4]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[4]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[4]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[4]_inst_i_5_n_0 ),
        .O(RD2_OBUF[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_10 
       (.I0(\r11_reg_n_0_[4] ),
        .I1(\r10_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_11 
       (.I0(\r15_reg_n_0_[4] ),
        .I1(\r14_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[4]_inst_i_12 
       (.I0(\r3_reg_n_0_[4] ),
        .I1(\r2_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_13 
       (.I0(\r7_reg_n_0_[4] ),
        .I1(\r6_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[4]_inst_i_2 
       (.I0(\RD2_OBUF[4]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[4]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[4]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[4]_inst_i_3 
       (.I0(\RD2_OBUF[4]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[4]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[4]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[4]_inst_i_4 
       (.I0(\RD2_OBUF[4]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[4]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[4]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[4]_inst_i_5 
       (.I0(\RD2_OBUF[4]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[4]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[4]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_6 
       (.I0(\r27_reg_n_0_[4] ),
        .I1(\r26_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_7 
       (.I0(\r31_reg_n_0_[4] ),
        .I1(\r30_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_8 
       (.I0(\r19_reg_n_0_[4] ),
        .I1(\r18_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[4]_inst_i_9 
       (.I0(\r23_reg_n_0_[4] ),
        .I1(\r22_reg_n_0_[4] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[4] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[4] ),
        .O(\RD2_OBUF[4]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[5]_inst 
       (.I(RD2_OBUF[5]),
        .O(RD2[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_1 
       (.I0(\RD2_OBUF[5]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[5]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[5]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[5]_inst_i_5_n_0 ),
        .O(RD2_OBUF[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_10 
       (.I0(\r11_reg_n_0_[5] ),
        .I1(\r10_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_11 
       (.I0(\r15_reg_n_0_[5] ),
        .I1(\r14_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[5]_inst_i_12 
       (.I0(\r3_reg_n_0_[5] ),
        .I1(\r2_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_13 
       (.I0(\r7_reg_n_0_[5] ),
        .I1(\r6_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[5]_inst_i_2 
       (.I0(\RD2_OBUF[5]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[5]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[5]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[5]_inst_i_3 
       (.I0(\RD2_OBUF[5]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[5]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[5]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[5]_inst_i_4 
       (.I0(\RD2_OBUF[5]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[5]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[5]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[5]_inst_i_5 
       (.I0(\RD2_OBUF[5]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[5]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[5]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_6 
       (.I0(\r27_reg_n_0_[5] ),
        .I1(\r26_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_7 
       (.I0(\r31_reg_n_0_[5] ),
        .I1(\r30_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_8 
       (.I0(\r19_reg_n_0_[5] ),
        .I1(\r18_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[5]_inst_i_9 
       (.I0(\r23_reg_n_0_[5] ),
        .I1(\r22_reg_n_0_[5] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[5] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[5] ),
        .O(\RD2_OBUF[5]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[6]_inst 
       (.I(RD2_OBUF[6]),
        .O(RD2[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_1 
       (.I0(\RD2_OBUF[6]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[6]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[6]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[6]_inst_i_5_n_0 ),
        .O(RD2_OBUF[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_10 
       (.I0(\r11_reg_n_0_[6] ),
        .I1(\r10_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_11 
       (.I0(\r15_reg_n_0_[6] ),
        .I1(\r14_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[6]_inst_i_12 
       (.I0(\r3_reg_n_0_[6] ),
        .I1(\r2_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_13 
       (.I0(\r7_reg_n_0_[6] ),
        .I1(\r6_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[6]_inst_i_2 
       (.I0(\RD2_OBUF[6]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[6]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[6]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[6]_inst_i_3 
       (.I0(\RD2_OBUF[6]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[6]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[6]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[6]_inst_i_4 
       (.I0(\RD2_OBUF[6]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[6]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[6]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[6]_inst_i_5 
       (.I0(\RD2_OBUF[6]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[6]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[6]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_6 
       (.I0(\r27_reg_n_0_[6] ),
        .I1(\r26_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_7 
       (.I0(\r31_reg_n_0_[6] ),
        .I1(\r30_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_8 
       (.I0(\r19_reg_n_0_[6] ),
        .I1(\r18_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[6]_inst_i_9 
       (.I0(\r23_reg_n_0_[6] ),
        .I1(\r22_reg_n_0_[6] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[6] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[6] ),
        .O(\RD2_OBUF[6]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[7]_inst 
       (.I(RD2_OBUF[7]),
        .O(RD2[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_1 
       (.I0(\RD2_OBUF[7]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[7]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[7]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[7]_inst_i_5_n_0 ),
        .O(RD2_OBUF[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_10 
       (.I0(\r11_reg_n_0_[7] ),
        .I1(\r10_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_11 
       (.I0(\r15_reg_n_0_[7] ),
        .I1(\r14_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[7]_inst_i_12 
       (.I0(\r3_reg_n_0_[7] ),
        .I1(\r2_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_13 
       (.I0(\r7_reg_n_0_[7] ),
        .I1(\r6_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[7]_inst_i_2 
       (.I0(\RD2_OBUF[7]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[7]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[7]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[7]_inst_i_3 
       (.I0(\RD2_OBUF[7]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[7]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[7]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[7]_inst_i_4 
       (.I0(\RD2_OBUF[7]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[7]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[7]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[7]_inst_i_5 
       (.I0(\RD2_OBUF[7]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[7]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[7]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_6 
       (.I0(\r27_reg_n_0_[7] ),
        .I1(\r26_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_7 
       (.I0(\r31_reg_n_0_[7] ),
        .I1(\r30_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_8 
       (.I0(\r19_reg_n_0_[7] ),
        .I1(\r18_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[7]_inst_i_9 
       (.I0(\r23_reg_n_0_[7] ),
        .I1(\r22_reg_n_0_[7] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[7] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[7] ),
        .O(\RD2_OBUF[7]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[8]_inst 
       (.I(RD2_OBUF[8]),
        .O(RD2[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_1 
       (.I0(\RD2_OBUF[8]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[8]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[8]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[8]_inst_i_5_n_0 ),
        .O(RD2_OBUF[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_10 
       (.I0(\r11_reg_n_0_[8] ),
        .I1(\r10_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_11 
       (.I0(\r15_reg_n_0_[8] ),
        .I1(\r14_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[8]_inst_i_12 
       (.I0(\r3_reg_n_0_[8] ),
        .I1(\r2_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_13 
       (.I0(\r7_reg_n_0_[8] ),
        .I1(\r6_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[8]_inst_i_2 
       (.I0(\RD2_OBUF[8]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[8]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[8]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[8]_inst_i_3 
       (.I0(\RD2_OBUF[8]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[8]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[8]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[8]_inst_i_4 
       (.I0(\RD2_OBUF[8]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[8]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[8]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[8]_inst_i_5 
       (.I0(\RD2_OBUF[8]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[8]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[8]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_6 
       (.I0(\r27_reg_n_0_[8] ),
        .I1(\r26_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_7 
       (.I0(\r31_reg_n_0_[8] ),
        .I1(\r30_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_8 
       (.I0(\r19_reg_n_0_[8] ),
        .I1(\r18_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[8]_inst_i_9 
       (.I0(\r23_reg_n_0_[8] ),
        .I1(\r22_reg_n_0_[8] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[8] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[8] ),
        .O(\RD2_OBUF[8]_inst_i_9_n_0 ));
  OBUF \RD2_OBUF[9]_inst 
       (.I(RD2_OBUF[9]),
        .O(RD2[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_1 
       (.I0(\RD2_OBUF[9]_inst_i_2_n_0 ),
        .I1(\RD2_OBUF[9]_inst_i_3_n_0 ),
        .I2(A2_IBUF[4]),
        .I3(\RD2_OBUF[9]_inst_i_4_n_0 ),
        .I4(A2_IBUF[3]),
        .I5(\RD2_OBUF[9]_inst_i_5_n_0 ),
        .O(RD2_OBUF[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_10 
       (.I0(\r11_reg_n_0_[9] ),
        .I1(\r10_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r9_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r8_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_11 
       (.I0(\r15_reg_n_0_[9] ),
        .I1(\r14_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r13_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r12_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \RD2_OBUF[9]_inst_i_12 
       (.I0(\r3_reg_n_0_[9] ),
        .I1(\r2_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(A2_IBUF[0]),
        .I4(\r1_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_13 
       (.I0(\r7_reg_n_0_[9] ),
        .I1(\r6_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r5_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r4_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_13_n_0 ));
  MUXF7 \RD2_OBUF[9]_inst_i_2 
       (.I0(\RD2_OBUF[9]_inst_i_6_n_0 ),
        .I1(\RD2_OBUF[9]_inst_i_7_n_0 ),
        .O(\RD2_OBUF[9]_inst_i_2_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[9]_inst_i_3 
       (.I0(\RD2_OBUF[9]_inst_i_8_n_0 ),
        .I1(\RD2_OBUF[9]_inst_i_9_n_0 ),
        .O(\RD2_OBUF[9]_inst_i_3_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[9]_inst_i_4 
       (.I0(\RD2_OBUF[9]_inst_i_10_n_0 ),
        .I1(\RD2_OBUF[9]_inst_i_11_n_0 ),
        .O(\RD2_OBUF[9]_inst_i_4_n_0 ),
        .S(A2_IBUF[2]));
  MUXF7 \RD2_OBUF[9]_inst_i_5 
       (.I0(\RD2_OBUF[9]_inst_i_12_n_0 ),
        .I1(\RD2_OBUF[9]_inst_i_13_n_0 ),
        .O(\RD2_OBUF[9]_inst_i_5_n_0 ),
        .S(A2_IBUF[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_6 
       (.I0(\r27_reg_n_0_[9] ),
        .I1(\r26_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r25_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r24_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_7 
       (.I0(\r31_reg_n_0_[9] ),
        .I1(\r30_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r29_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r28_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_8 
       (.I0(\r19_reg_n_0_[9] ),
        .I1(\r18_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r17_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r16_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \RD2_OBUF[9]_inst_i_9 
       (.I0(\r23_reg_n_0_[9] ),
        .I1(\r22_reg_n_0_[9] ),
        .I2(A2_IBUF[1]),
        .I3(\r21_reg_n_0_[9] ),
        .I4(A2_IBUF[0]),
        .I5(\r20_reg_n_0_[9] ),
        .O(\RD2_OBUF[9]_inst_i_9_n_0 ));
  IBUF \WD_IBUF[0]_inst 
       (.I(WD[0]),
        .O(WD_IBUF[0]));
  IBUF \WD_IBUF[10]_inst 
       (.I(WD[10]),
        .O(WD_IBUF[10]));
  IBUF \WD_IBUF[11]_inst 
       (.I(WD[11]),
        .O(WD_IBUF[11]));
  IBUF \WD_IBUF[12]_inst 
       (.I(WD[12]),
        .O(WD_IBUF[12]));
  IBUF \WD_IBUF[13]_inst 
       (.I(WD[13]),
        .O(WD_IBUF[13]));
  IBUF \WD_IBUF[14]_inst 
       (.I(WD[14]),
        .O(WD_IBUF[14]));
  IBUF \WD_IBUF[15]_inst 
       (.I(WD[15]),
        .O(WD_IBUF[15]));
  IBUF \WD_IBUF[16]_inst 
       (.I(WD[16]),
        .O(WD_IBUF[16]));
  IBUF \WD_IBUF[17]_inst 
       (.I(WD[17]),
        .O(WD_IBUF[17]));
  IBUF \WD_IBUF[18]_inst 
       (.I(WD[18]),
        .O(WD_IBUF[18]));
  IBUF \WD_IBUF[19]_inst 
       (.I(WD[19]),
        .O(WD_IBUF[19]));
  IBUF \WD_IBUF[1]_inst 
       (.I(WD[1]),
        .O(WD_IBUF[1]));
  IBUF \WD_IBUF[20]_inst 
       (.I(WD[20]),
        .O(WD_IBUF[20]));
  IBUF \WD_IBUF[21]_inst 
       (.I(WD[21]),
        .O(WD_IBUF[21]));
  IBUF \WD_IBUF[22]_inst 
       (.I(WD[22]),
        .O(WD_IBUF[22]));
  IBUF \WD_IBUF[23]_inst 
       (.I(WD[23]),
        .O(WD_IBUF[23]));
  IBUF \WD_IBUF[24]_inst 
       (.I(WD[24]),
        .O(WD_IBUF[24]));
  IBUF \WD_IBUF[25]_inst 
       (.I(WD[25]),
        .O(WD_IBUF[25]));
  IBUF \WD_IBUF[26]_inst 
       (.I(WD[26]),
        .O(WD_IBUF[26]));
  IBUF \WD_IBUF[27]_inst 
       (.I(WD[27]),
        .O(WD_IBUF[27]));
  IBUF \WD_IBUF[28]_inst 
       (.I(WD[28]),
        .O(WD_IBUF[28]));
  IBUF \WD_IBUF[29]_inst 
       (.I(WD[29]),
        .O(WD_IBUF[29]));
  IBUF \WD_IBUF[2]_inst 
       (.I(WD[2]),
        .O(WD_IBUF[2]));
  IBUF \WD_IBUF[30]_inst 
       (.I(WD[30]),
        .O(WD_IBUF[30]));
  IBUF \WD_IBUF[31]_inst 
       (.I(WD[31]),
        .O(WD_IBUF[31]));
  IBUF \WD_IBUF[3]_inst 
       (.I(WD[3]),
        .O(WD_IBUF[3]));
  IBUF \WD_IBUF[4]_inst 
       (.I(WD[4]),
        .O(WD_IBUF[4]));
  IBUF \WD_IBUF[5]_inst 
       (.I(WD[5]),
        .O(WD_IBUF[5]));
  IBUF \WD_IBUF[6]_inst 
       (.I(WD[6]),
        .O(WD_IBUF[6]));
  IBUF \WD_IBUF[7]_inst 
       (.I(WD[7]),
        .O(WD_IBUF[7]));
  IBUF \WD_IBUF[8]_inst 
       (.I(WD[8]),
        .O(WD_IBUF[8]));
  IBUF \WD_IBUF[9]_inst 
       (.I(WD[9]),
        .O(WD_IBUF[9]));
  IBUF WE_IBUF_inst
       (.I(WE),
        .O(WE_IBUF));
  BUFG clk_IBUF_BUFG_inst
       (.I(clk_IBUF),
        .O(clk_IBUF_BUFG));
  IBUF clk_IBUF_inst
       (.I(clk),
        .O(clk_IBUF));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r10[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[2]),
        .O(r10));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[0]),
        .Q(\r10_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[10]),
        .Q(\r10_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[11]),
        .Q(\r10_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[12]),
        .Q(\r10_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[13]),
        .Q(\r10_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[14]),
        .Q(\r10_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[15]),
        .Q(\r10_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[16]),
        .Q(\r10_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[17]),
        .Q(\r10_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[18]),
        .Q(\r10_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[19]),
        .Q(\r10_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[1]),
        .Q(\r10_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[20]),
        .Q(\r10_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[21]),
        .Q(\r10_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[22]),
        .Q(\r10_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[23]),
        .Q(\r10_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[24]),
        .Q(\r10_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[25]),
        .Q(\r10_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[26]),
        .Q(\r10_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[27]),
        .Q(\r10_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[28]),
        .Q(\r10_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[29]),
        .Q(\r10_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[2]),
        .Q(\r10_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[30]),
        .Q(\r10_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[31]),
        .Q(\r10_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[3]),
        .Q(\r10_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[4]),
        .Q(\r10_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[5]),
        .Q(\r10_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[6]),
        .Q(\r10_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[7]),
        .Q(\r10_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[8]),
        .Q(\r10_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r10_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r10),
        .D(WD_IBUF[9]),
        .Q(\r10_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r11[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[2]),
        .O(r11));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[0]),
        .Q(\r11_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[10]),
        .Q(\r11_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[11]),
        .Q(\r11_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[12]),
        .Q(\r11_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[13]),
        .Q(\r11_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[14]),
        .Q(\r11_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[15]),
        .Q(\r11_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[16]),
        .Q(\r11_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[17]),
        .Q(\r11_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[18]),
        .Q(\r11_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[19]),
        .Q(\r11_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[1]),
        .Q(\r11_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[20]),
        .Q(\r11_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[21]),
        .Q(\r11_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[22]),
        .Q(\r11_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[23]),
        .Q(\r11_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[24]),
        .Q(\r11_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[25]),
        .Q(\r11_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[26]),
        .Q(\r11_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[27]),
        .Q(\r11_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[28]),
        .Q(\r11_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[29]),
        .Q(\r11_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[2]),
        .Q(\r11_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[30]),
        .Q(\r11_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[31]),
        .Q(\r11_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[3]),
        .Q(\r11_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[4]),
        .Q(\r11_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[5]),
        .Q(\r11_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[6]),
        .Q(\r11_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[7]),
        .Q(\r11_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[8]),
        .Q(\r11_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r11_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r11),
        .D(WD_IBUF[9]),
        .Q(\r11_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r12[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[1]),
        .O(r12));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[0]),
        .Q(\r12_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[10]),
        .Q(\r12_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[11]),
        .Q(\r12_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[12]),
        .Q(\r12_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[13]),
        .Q(\r12_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[14]),
        .Q(\r12_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[15]),
        .Q(\r12_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[16]),
        .Q(\r12_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[17]),
        .Q(\r12_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[18]),
        .Q(\r12_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[19]),
        .Q(\r12_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[1]),
        .Q(\r12_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[20]),
        .Q(\r12_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[21]),
        .Q(\r12_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[22]),
        .Q(\r12_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[23]),
        .Q(\r12_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[24]),
        .Q(\r12_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[25]),
        .Q(\r12_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[26]),
        .Q(\r12_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[27]),
        .Q(\r12_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[28]),
        .Q(\r12_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[29]),
        .Q(\r12_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[2]),
        .Q(\r12_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[30]),
        .Q(\r12_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[31]),
        .Q(\r12_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[3]),
        .Q(\r12_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[4]),
        .Q(\r12_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[5]),
        .Q(\r12_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[6]),
        .Q(\r12_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[7]),
        .Q(\r12_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[8]),
        .Q(\r12_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r12_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r12),
        .D(WD_IBUF[9]),
        .Q(\r12_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r13[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[1]),
        .O(r13));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[0]),
        .Q(\r13_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[10]),
        .Q(\r13_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[11]),
        .Q(\r13_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[12]),
        .Q(\r13_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[13]),
        .Q(\r13_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[14]),
        .Q(\r13_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[15]),
        .Q(\r13_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[16]),
        .Q(\r13_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[17]),
        .Q(\r13_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[18]),
        .Q(\r13_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[19]),
        .Q(\r13_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[1]),
        .Q(\r13_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[20]),
        .Q(\r13_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[21]),
        .Q(\r13_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[22]),
        .Q(\r13_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[23]),
        .Q(\r13_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[24]),
        .Q(\r13_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[25]),
        .Q(\r13_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[26]),
        .Q(\r13_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[27]),
        .Q(\r13_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[28]),
        .Q(\r13_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[29]),
        .Q(\r13_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[2]),
        .Q(\r13_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[30]),
        .Q(\r13_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[31]),
        .Q(\r13_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[3]),
        .Q(\r13_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[4]),
        .Q(\r13_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[5]),
        .Q(\r13_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[6]),
        .Q(\r13_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[7]),
        .Q(\r13_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[8]),
        .Q(\r13_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r13_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r13),
        .D(WD_IBUF[9]),
        .Q(\r13_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r14[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[0]),
        .O(r14));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[0]),
        .Q(\r14_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[10]),
        .Q(\r14_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[11]),
        .Q(\r14_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[12]),
        .Q(\r14_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[13]),
        .Q(\r14_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[14]),
        .Q(\r14_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[15]),
        .Q(\r14_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[16]),
        .Q(\r14_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[17]),
        .Q(\r14_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[18]),
        .Q(\r14_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[19]),
        .Q(\r14_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[1]),
        .Q(\r14_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[20]),
        .Q(\r14_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[21]),
        .Q(\r14_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[22]),
        .Q(\r14_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[23]),
        .Q(\r14_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[24]),
        .Q(\r14_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[25]),
        .Q(\r14_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[26]),
        .Q(\r14_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[27]),
        .Q(\r14_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[28]),
        .Q(\r14_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[29]),
        .Q(\r14_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[2]),
        .Q(\r14_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[30]),
        .Q(\r14_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[31]),
        .Q(\r14_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[3]),
        .Q(\r14_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[4]),
        .Q(\r14_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[5]),
        .Q(\r14_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[6]),
        .Q(\r14_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[7]),
        .Q(\r14_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[8]),
        .Q(\r14_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r14_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r14),
        .D(WD_IBUF[9]),
        .Q(\r14_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r15[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[3]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[1]),
        .I5(A3_IBUF[2]),
        .O(r15));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[0]),
        .Q(\r15_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[10]),
        .Q(\r15_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[11]),
        .Q(\r15_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[12]),
        .Q(\r15_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[13]),
        .Q(\r15_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[14]),
        .Q(\r15_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[15]),
        .Q(\r15_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[16]),
        .Q(\r15_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[17]),
        .Q(\r15_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[18]),
        .Q(\r15_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[19]),
        .Q(\r15_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[1]),
        .Q(\r15_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[20]),
        .Q(\r15_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[21]),
        .Q(\r15_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[22]),
        .Q(\r15_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[23]),
        .Q(\r15_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[24]),
        .Q(\r15_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[25]),
        .Q(\r15_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[26]),
        .Q(\r15_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[27]),
        .Q(\r15_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[28]),
        .Q(\r15_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[29]),
        .Q(\r15_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[2]),
        .Q(\r15_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[30]),
        .Q(\r15_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[31]),
        .Q(\r15_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[3]),
        .Q(\r15_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[4]),
        .Q(\r15_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[5]),
        .Q(\r15_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[6]),
        .Q(\r15_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[7]),
        .Q(\r15_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[8]),
        .Q(\r15_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r15_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r15),
        .D(WD_IBUF[9]),
        .Q(\r15_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r16[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[4]),
        .I4(A3_IBUF[0]),
        .I5(A3_IBUF[2]),
        .O(r16));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[0]),
        .Q(\r16_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[10]),
        .Q(\r16_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[11]),
        .Q(\r16_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[12]),
        .Q(\r16_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[13]),
        .Q(\r16_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[14]),
        .Q(\r16_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[15]),
        .Q(\r16_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[16]),
        .Q(\r16_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[17]),
        .Q(\r16_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[18]),
        .Q(\r16_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[19]),
        .Q(\r16_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[1]),
        .Q(\r16_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[20]),
        .Q(\r16_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[21]),
        .Q(\r16_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[22]),
        .Q(\r16_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[23]),
        .Q(\r16_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[24]),
        .Q(\r16_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[25]),
        .Q(\r16_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[26]),
        .Q(\r16_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[27]),
        .Q(\r16_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[28]),
        .Q(\r16_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[29]),
        .Q(\r16_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[2]),
        .Q(\r16_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[30]),
        .Q(\r16_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[31]),
        .Q(\r16_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[3]),
        .Q(\r16_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[4]),
        .Q(\r16_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[5]),
        .Q(\r16_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[6]),
        .Q(\r16_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[7]),
        .Q(\r16_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[8]),
        .Q(\r16_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r16_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r16),
        .D(WD_IBUF[9]),
        .Q(\r16_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r17[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[2]),
        .O(r17));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[0]),
        .Q(\r17_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[10]),
        .Q(\r17_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[11]),
        .Q(\r17_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[12]),
        .Q(\r17_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[13]),
        .Q(\r17_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[14]),
        .Q(\r17_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[15]),
        .Q(\r17_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[16]),
        .Q(\r17_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[17]),
        .Q(\r17_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[18]),
        .Q(\r17_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[19]),
        .Q(\r17_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[1]),
        .Q(\r17_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[20]),
        .Q(\r17_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[21]),
        .Q(\r17_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[22]),
        .Q(\r17_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[23]),
        .Q(\r17_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[24]),
        .Q(\r17_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[25]),
        .Q(\r17_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[26]),
        .Q(\r17_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[27]),
        .Q(\r17_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[28]),
        .Q(\r17_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[29]),
        .Q(\r17_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[2]),
        .Q(\r17_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[30]),
        .Q(\r17_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[31]),
        .Q(\r17_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[3]),
        .Q(\r17_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[4]),
        .Q(\r17_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[5]),
        .Q(\r17_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[6]),
        .Q(\r17_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[7]),
        .Q(\r17_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[8]),
        .Q(\r17_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r17_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r17),
        .D(WD_IBUF[9]),
        .Q(\r17_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r18[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[2]),
        .O(r18));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[0]),
        .Q(\r18_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[10]),
        .Q(\r18_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[11]),
        .Q(\r18_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[12]),
        .Q(\r18_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[13]),
        .Q(\r18_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[14]),
        .Q(\r18_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[15]),
        .Q(\r18_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[16]),
        .Q(\r18_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[17]),
        .Q(\r18_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[18]),
        .Q(\r18_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[19]),
        .Q(\r18_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[1]),
        .Q(\r18_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[20]),
        .Q(\r18_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[21]),
        .Q(\r18_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[22]),
        .Q(\r18_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[23]),
        .Q(\r18_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[24]),
        .Q(\r18_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[25]),
        .Q(\r18_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[26]),
        .Q(\r18_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[27]),
        .Q(\r18_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[28]),
        .Q(\r18_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[29]),
        .Q(\r18_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[2]),
        .Q(\r18_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[30]),
        .Q(\r18_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[31]),
        .Q(\r18_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[3]),
        .Q(\r18_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[4]),
        .Q(\r18_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[5]),
        .Q(\r18_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[6]),
        .Q(\r18_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[7]),
        .Q(\r18_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[8]),
        .Q(\r18_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r18_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r18),
        .D(WD_IBUF[9]),
        .Q(\r18_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r19[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[2]),
        .O(r19));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[0]),
        .Q(\r19_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[10]),
        .Q(\r19_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[11]),
        .Q(\r19_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[12]),
        .Q(\r19_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[13]),
        .Q(\r19_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[14]),
        .Q(\r19_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[15]),
        .Q(\r19_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[16]),
        .Q(\r19_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[17]),
        .Q(\r19_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[18]),
        .Q(\r19_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[19]),
        .Q(\r19_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[1]),
        .Q(\r19_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[20]),
        .Q(\r19_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[21]),
        .Q(\r19_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[22]),
        .Q(\r19_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[23]),
        .Q(\r19_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[24]),
        .Q(\r19_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[25]),
        .Q(\r19_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[26]),
        .Q(\r19_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[27]),
        .Q(\r19_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[28]),
        .Q(\r19_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[29]),
        .Q(\r19_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[2]),
        .Q(\r19_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[30]),
        .Q(\r19_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[31]),
        .Q(\r19_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[3]),
        .Q(\r19_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[4]),
        .Q(\r19_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[5]),
        .Q(\r19_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[6]),
        .Q(\r19_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[7]),
        .Q(\r19_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[8]),
        .Q(\r19_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r19_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r19),
        .D(WD_IBUF[9]),
        .Q(\r19_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r1[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[2]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[1]),
        .I5(A3_IBUF[4]),
        .O(r1));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[0]),
        .Q(\r1_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[10]),
        .Q(\r1_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[11]),
        .Q(\r1_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[12]),
        .Q(\r1_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[13]),
        .Q(\r1_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[14]),
        .Q(\r1_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[15]),
        .Q(\r1_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[16]),
        .Q(\r1_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[17]),
        .Q(\r1_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[18]),
        .Q(\r1_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[19]),
        .Q(\r1_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[1]),
        .Q(\r1_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[20]),
        .Q(\r1_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[21]),
        .Q(\r1_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[22]),
        .Q(\r1_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[23]),
        .Q(\r1_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[24]),
        .Q(\r1_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[25]),
        .Q(\r1_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[26]),
        .Q(\r1_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[27]),
        .Q(\r1_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[28]),
        .Q(\r1_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[29]),
        .Q(\r1_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[2]),
        .Q(\r1_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[30]),
        .Q(\r1_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[31]),
        .Q(\r1_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[3]),
        .Q(\r1_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[4]),
        .Q(\r1_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[5]),
        .Q(\r1_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[6]),
        .Q(\r1_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[7]),
        .Q(\r1_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[8]),
        .Q(\r1_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r1_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r1),
        .D(WD_IBUF[9]),
        .Q(\r1_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r20[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[1]),
        .O(r20));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[0]),
        .Q(\r20_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[10]),
        .Q(\r20_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[11]),
        .Q(\r20_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[12]),
        .Q(\r20_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[13]),
        .Q(\r20_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[14]),
        .Q(\r20_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[15]),
        .Q(\r20_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[16]),
        .Q(\r20_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[17]),
        .Q(\r20_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[18]),
        .Q(\r20_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[19]),
        .Q(\r20_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[1]),
        .Q(\r20_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[20]),
        .Q(\r20_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[21]),
        .Q(\r20_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[22]),
        .Q(\r20_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[23]),
        .Q(\r20_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[24]),
        .Q(\r20_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[25]),
        .Q(\r20_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[26]),
        .Q(\r20_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[27]),
        .Q(\r20_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[28]),
        .Q(\r20_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[29]),
        .Q(\r20_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[2]),
        .Q(\r20_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[30]),
        .Q(\r20_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[31]),
        .Q(\r20_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[3]),
        .Q(\r20_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[4]),
        .Q(\r20_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[5]),
        .Q(\r20_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[6]),
        .Q(\r20_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[7]),
        .Q(\r20_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[8]),
        .Q(\r20_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r20_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r20),
        .D(WD_IBUF[9]),
        .Q(\r20_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r21[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[1]),
        .O(r21));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[0]),
        .Q(\r21_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[10]),
        .Q(\r21_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[11]),
        .Q(\r21_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[12]),
        .Q(\r21_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[13]),
        .Q(\r21_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[14]),
        .Q(\r21_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[15]),
        .Q(\r21_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[16]),
        .Q(\r21_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[17]),
        .Q(\r21_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[18]),
        .Q(\r21_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[19]),
        .Q(\r21_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[1]),
        .Q(\r21_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[20]),
        .Q(\r21_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[21]),
        .Q(\r21_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[22]),
        .Q(\r21_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[23]),
        .Q(\r21_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[24]),
        .Q(\r21_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[25]),
        .Q(\r21_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[26]),
        .Q(\r21_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[27]),
        .Q(\r21_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[28]),
        .Q(\r21_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[29]),
        .Q(\r21_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[2]),
        .Q(\r21_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[30]),
        .Q(\r21_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[31]),
        .Q(\r21_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[3]),
        .Q(\r21_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[4]),
        .Q(\r21_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[5]),
        .Q(\r21_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[6]),
        .Q(\r21_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[7]),
        .Q(\r21_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[8]),
        .Q(\r21_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r21_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r21),
        .D(WD_IBUF[9]),
        .Q(\r21_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r22[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[0]),
        .O(r22));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[0]),
        .Q(\r22_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[10]),
        .Q(\r22_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[11]),
        .Q(\r22_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[12]),
        .Q(\r22_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[13]),
        .Q(\r22_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[14]),
        .Q(\r22_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[15]),
        .Q(\r22_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[16]),
        .Q(\r22_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[17]),
        .Q(\r22_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[18]),
        .Q(\r22_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[19]),
        .Q(\r22_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[1]),
        .Q(\r22_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[20]),
        .Q(\r22_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[21]),
        .Q(\r22_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[22]),
        .Q(\r22_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[23]),
        .Q(\r22_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[24]),
        .Q(\r22_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[25]),
        .Q(\r22_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[26]),
        .Q(\r22_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[27]),
        .Q(\r22_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[28]),
        .Q(\r22_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[29]),
        .Q(\r22_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[2]),
        .Q(\r22_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[30]),
        .Q(\r22_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[31]),
        .Q(\r22_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[3]),
        .Q(\r22_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[4]),
        .Q(\r22_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[5]),
        .Q(\r22_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[6]),
        .Q(\r22_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[7]),
        .Q(\r22_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[8]),
        .Q(\r22_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r22_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r22),
        .D(WD_IBUF[9]),
        .Q(\r22_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r23[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[4]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[1]),
        .I5(A3_IBUF[2]),
        .O(r23));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[0]),
        .Q(\r23_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[10]),
        .Q(\r23_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[11]),
        .Q(\r23_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[12]),
        .Q(\r23_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[13]),
        .Q(\r23_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[14]),
        .Q(\r23_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[15]),
        .Q(\r23_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[16]),
        .Q(\r23_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[17]),
        .Q(\r23_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[18]),
        .Q(\r23_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[19]),
        .Q(\r23_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[1]),
        .Q(\r23_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[20]),
        .Q(\r23_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[21]),
        .Q(\r23_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[22]),
        .Q(\r23_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[23]),
        .Q(\r23_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[24]),
        .Q(\r23_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[25]),
        .Q(\r23_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[26]),
        .Q(\r23_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[27]),
        .Q(\r23_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[28]),
        .Q(\r23_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[29]),
        .Q(\r23_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[2]),
        .Q(\r23_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[30]),
        .Q(\r23_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[31]),
        .Q(\r23_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[3]),
        .Q(\r23_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[4]),
        .Q(\r23_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[5]),
        .Q(\r23_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[6]),
        .Q(\r23_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[7]),
        .Q(\r23_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[8]),
        .Q(\r23_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r23_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r23),
        .D(WD_IBUF[9]),
        .Q(\r23_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r24[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[2]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[4]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[1]),
        .O(r24));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[0]),
        .Q(\r24_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[10]),
        .Q(\r24_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[11]),
        .Q(\r24_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[12]),
        .Q(\r24_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[13]),
        .Q(\r24_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[14]),
        .Q(\r24_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[15]),
        .Q(\r24_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[16]),
        .Q(\r24_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[17]),
        .Q(\r24_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[18]),
        .Q(\r24_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[19]),
        .Q(\r24_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[1]),
        .Q(\r24_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[20]),
        .Q(\r24_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[21]),
        .Q(\r24_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[22]),
        .Q(\r24_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[23]),
        .Q(\r24_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[24]),
        .Q(\r24_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[25]),
        .Q(\r24_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[26]),
        .Q(\r24_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[27]),
        .Q(\r24_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[28]),
        .Q(\r24_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[29]),
        .Q(\r24_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[2]),
        .Q(\r24_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[30]),
        .Q(\r24_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[31]),
        .Q(\r24_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[3]),
        .Q(\r24_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[4]),
        .Q(\r24_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[5]),
        .Q(\r24_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[6]),
        .Q(\r24_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[7]),
        .Q(\r24_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[8]),
        .Q(\r24_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r24_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r24),
        .D(WD_IBUF[9]),
        .Q(\r24_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r25[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[2]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[4]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[1]),
        .O(r25));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[0]),
        .Q(\r25_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[10]),
        .Q(\r25_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[11]),
        .Q(\r25_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[12]),
        .Q(\r25_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[13]),
        .Q(\r25_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[14]),
        .Q(\r25_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[15]),
        .Q(\r25_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[16]),
        .Q(\r25_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[17]),
        .Q(\r25_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[18]),
        .Q(\r25_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[19]),
        .Q(\r25_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[1]),
        .Q(\r25_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[20]),
        .Q(\r25_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[21]),
        .Q(\r25_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[22]),
        .Q(\r25_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[23]),
        .Q(\r25_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[24]),
        .Q(\r25_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[25]),
        .Q(\r25_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[26]),
        .Q(\r25_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[27]),
        .Q(\r25_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[28]),
        .Q(\r25_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[29]),
        .Q(\r25_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[2]),
        .Q(\r25_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[30]),
        .Q(\r25_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[31]),
        .Q(\r25_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[3]),
        .Q(\r25_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[4]),
        .Q(\r25_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[5]),
        .Q(\r25_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[6]),
        .Q(\r25_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[7]),
        .Q(\r25_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[8]),
        .Q(\r25_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r25_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r25),
        .D(WD_IBUF[9]),
        .Q(\r25_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r26[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[2]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[4]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[0]),
        .O(r26));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[0]),
        .Q(\r26_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[10]),
        .Q(\r26_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[11]),
        .Q(\r26_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[12]),
        .Q(\r26_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[13]),
        .Q(\r26_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[14]),
        .Q(\r26_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[15]),
        .Q(\r26_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[16]),
        .Q(\r26_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[17]),
        .Q(\r26_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[18]),
        .Q(\r26_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[19]),
        .Q(\r26_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[1]),
        .Q(\r26_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[20]),
        .Q(\r26_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[21]),
        .Q(\r26_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[22]),
        .Q(\r26_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[23]),
        .Q(\r26_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[24]),
        .Q(\r26_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[25]),
        .Q(\r26_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[26]),
        .Q(\r26_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[27]),
        .Q(\r26_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[28]),
        .Q(\r26_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[29]),
        .Q(\r26_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[2]),
        .Q(\r26_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[30]),
        .Q(\r26_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[31]),
        .Q(\r26_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[3]),
        .Q(\r26_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[4]),
        .Q(\r26_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[5]),
        .Q(\r26_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[6]),
        .Q(\r26_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[7]),
        .Q(\r26_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[8]),
        .Q(\r26_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r26_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r26),
        .D(WD_IBUF[9]),
        .Q(\r26_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r27[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[2]),
        .I2(A3_IBUF[3]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[1]),
        .I5(A3_IBUF[4]),
        .O(r27));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[0]),
        .Q(\r27_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[10]),
        .Q(\r27_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[11]),
        .Q(\r27_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[12]),
        .Q(\r27_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[13]),
        .Q(\r27_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[14]),
        .Q(\r27_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[15]),
        .Q(\r27_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[16]),
        .Q(\r27_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[17]),
        .Q(\r27_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[18]),
        .Q(\r27_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[19]),
        .Q(\r27_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[1]),
        .Q(\r27_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[20]),
        .Q(\r27_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[21]),
        .Q(\r27_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[22]),
        .Q(\r27_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[23]),
        .Q(\r27_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[24]),
        .Q(\r27_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[25]),
        .Q(\r27_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[26]),
        .Q(\r27_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[27]),
        .Q(\r27_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[28]),
        .Q(\r27_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[29]),
        .Q(\r27_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[2]),
        .Q(\r27_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[30]),
        .Q(\r27_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[31]),
        .Q(\r27_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[3]),
        .Q(\r27_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[4]),
        .Q(\r27_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[5]),
        .Q(\r27_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[6]),
        .Q(\r27_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[7]),
        .Q(\r27_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[8]),
        .Q(\r27_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r27_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r27),
        .D(WD_IBUF[9]),
        .Q(\r27_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r28[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[1]),
        .I2(A3_IBUF[2]),
        .I3(A3_IBUF[4]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[0]),
        .O(r28));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[0]),
        .Q(\r28_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[10]),
        .Q(\r28_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[11]),
        .Q(\r28_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[12]),
        .Q(\r28_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[13]),
        .Q(\r28_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[14]),
        .Q(\r28_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[15]),
        .Q(\r28_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[16]),
        .Q(\r28_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[17]),
        .Q(\r28_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[18]),
        .Q(\r28_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[19]),
        .Q(\r28_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[1]),
        .Q(\r28_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[20]),
        .Q(\r28_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[21]),
        .Q(\r28_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[22]),
        .Q(\r28_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[23]),
        .Q(\r28_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[24]),
        .Q(\r28_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[25]),
        .Q(\r28_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[26]),
        .Q(\r28_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[27]),
        .Q(\r28_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[28]),
        .Q(\r28_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[29]),
        .Q(\r28_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[2]),
        .Q(\r28_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[30]),
        .Q(\r28_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[31]),
        .Q(\r28_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[3]),
        .Q(\r28_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[4]),
        .Q(\r28_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[5]),
        .Q(\r28_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[6]),
        .Q(\r28_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[7]),
        .Q(\r28_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[8]),
        .Q(\r28_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r28_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r28),
        .D(WD_IBUF[9]),
        .Q(\r28_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r29[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[1]),
        .I2(A3_IBUF[3]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[2]),
        .I5(A3_IBUF[4]),
        .O(r29));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[0]),
        .Q(\r29_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[10]),
        .Q(\r29_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[11]),
        .Q(\r29_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[12]),
        .Q(\r29_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[13]),
        .Q(\r29_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[14]),
        .Q(\r29_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[15]),
        .Q(\r29_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[16]),
        .Q(\r29_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[17]),
        .Q(\r29_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[18]),
        .Q(\r29_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[19]),
        .Q(\r29_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[1]),
        .Q(\r29_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[20]),
        .Q(\r29_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[21]),
        .Q(\r29_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[22]),
        .Q(\r29_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[23]),
        .Q(\r29_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[24]),
        .Q(\r29_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[25]),
        .Q(\r29_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[26]),
        .Q(\r29_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[27]),
        .Q(\r29_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[28]),
        .Q(\r29_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[29]),
        .Q(\r29_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[2]),
        .Q(\r29_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[30]),
        .Q(\r29_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[31]),
        .Q(\r29_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[3]),
        .Q(\r29_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[4]),
        .Q(\r29_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[5]),
        .Q(\r29_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[6]),
        .Q(\r29_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[7]),
        .Q(\r29_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[8]),
        .Q(\r29_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r29_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r29),
        .D(WD_IBUF[9]),
        .Q(\r29_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r2[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[2]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[0]),
        .I5(A3_IBUF[4]),
        .O(r2));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[0]),
        .Q(\r2_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[10]),
        .Q(\r2_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[11]),
        .Q(\r2_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[12]),
        .Q(\r2_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[13]),
        .Q(\r2_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[14]),
        .Q(\r2_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[15]),
        .Q(\r2_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[16]),
        .Q(\r2_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[17]),
        .Q(\r2_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[18]),
        .Q(\r2_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[19]),
        .Q(\r2_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[1]),
        .Q(\r2_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[20]),
        .Q(\r2_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[21]),
        .Q(\r2_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[22]),
        .Q(\r2_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[23]),
        .Q(\r2_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[24]),
        .Q(\r2_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[25]),
        .Q(\r2_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[26]),
        .Q(\r2_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[27]),
        .Q(\r2_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[28]),
        .Q(\r2_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[29]),
        .Q(\r2_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[2]),
        .Q(\r2_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[30]),
        .Q(\r2_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[31]),
        .Q(\r2_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[3]),
        .Q(\r2_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[4]),
        .Q(\r2_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[5]),
        .Q(\r2_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[6]),
        .Q(\r2_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[7]),
        .Q(\r2_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[8]),
        .Q(\r2_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r2_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r2),
        .D(WD_IBUF[9]),
        .Q(\r2_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r30[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[0]),
        .I2(A3_IBUF[3]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[2]),
        .I5(A3_IBUF[4]),
        .O(r30));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[0]),
        .Q(\r30_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[10]),
        .Q(\r30_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[11]),
        .Q(\r30_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[12]),
        .Q(\r30_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[13]),
        .Q(\r30_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[14]),
        .Q(\r30_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[15]),
        .Q(\r30_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[16]),
        .Q(\r30_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[17]),
        .Q(\r30_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[18]),
        .Q(\r30_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[19]),
        .Q(\r30_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[1]),
        .Q(\r30_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[20]),
        .Q(\r30_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[21]),
        .Q(\r30_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[22]),
        .Q(\r30_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[23]),
        .Q(\r30_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[24]),
        .Q(\r30_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[25]),
        .Q(\r30_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[26]),
        .Q(\r30_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[27]),
        .Q(\r30_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[28]),
        .Q(\r30_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[29]),
        .Q(\r30_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[2]),
        .Q(\r30_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[30]),
        .Q(\r30_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[31]),
        .Q(\r30_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[3]),
        .Q(\r30_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[4]),
        .Q(\r30_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[5]),
        .Q(\r30_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[6]),
        .Q(\r30_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[7]),
        .Q(\r30_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[8]),
        .Q(\r30_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r30_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r30),
        .D(WD_IBUF[9]),
        .Q(\r30_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r31[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[2]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[4]),
        .I5(A3_IBUF[3]),
        .O(r31));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[0]),
        .Q(\r31_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[10]),
        .Q(\r31_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[11]),
        .Q(\r31_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[12]),
        .Q(\r31_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[13]),
        .Q(\r31_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[14]),
        .Q(\r31_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[15]),
        .Q(\r31_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[16]),
        .Q(\r31_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[17]),
        .Q(\r31_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[18]),
        .Q(\r31_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[19]),
        .Q(\r31_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[1]),
        .Q(\r31_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[20]),
        .Q(\r31_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[21]),
        .Q(\r31_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[22]),
        .Q(\r31_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[23]),
        .Q(\r31_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[24]),
        .Q(\r31_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[25]),
        .Q(\r31_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[26]),
        .Q(\r31_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[27]),
        .Q(\r31_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[28]),
        .Q(\r31_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[29]),
        .Q(\r31_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[2]),
        .Q(\r31_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[30]),
        .Q(\r31_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[31]),
        .Q(\r31_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[3]),
        .Q(\r31_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[4]),
        .Q(\r31_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[5]),
        .Q(\r31_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[6]),
        .Q(\r31_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[7]),
        .Q(\r31_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[8]),
        .Q(\r31_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r31_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r31),
        .D(WD_IBUF[9]),
        .Q(\r31_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r3[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[2]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[1]),
        .I5(A3_IBUF[4]),
        .O(r3));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[0]),
        .Q(\r3_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[10]),
        .Q(\r3_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[11]),
        .Q(\r3_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[12]),
        .Q(\r3_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[13]),
        .Q(\r3_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[14]),
        .Q(\r3_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[15]),
        .Q(\r3_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[16]),
        .Q(\r3_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[17]),
        .Q(\r3_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[18]),
        .Q(\r3_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[19]),
        .Q(\r3_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[1]),
        .Q(\r3_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[20]),
        .Q(\r3_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[21]),
        .Q(\r3_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[22]),
        .Q(\r3_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[23]),
        .Q(\r3_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[24]),
        .Q(\r3_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[25]),
        .Q(\r3_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[26]),
        .Q(\r3_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[27]),
        .Q(\r3_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[28]),
        .Q(\r3_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[29]),
        .Q(\r3_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[2]),
        .Q(\r3_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[30]),
        .Q(\r3_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[31]),
        .Q(\r3_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[3]),
        .Q(\r3_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[4]),
        .Q(\r3_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[5]),
        .Q(\r3_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[6]),
        .Q(\r3_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[7]),
        .Q(\r3_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[8]),
        .Q(\r3_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r3_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r3),
        .D(WD_IBUF[9]),
        .Q(\r3_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r4[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[2]),
        .I4(A3_IBUF[0]),
        .I5(A3_IBUF[4]),
        .O(r4));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[0]),
        .Q(\r4_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[10]),
        .Q(\r4_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[11]),
        .Q(\r4_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[12]),
        .Q(\r4_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[13]),
        .Q(\r4_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[14]),
        .Q(\r4_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[15]),
        .Q(\r4_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[16]),
        .Q(\r4_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[17]),
        .Q(\r4_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[18]),
        .Q(\r4_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[19]),
        .Q(\r4_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[1]),
        .Q(\r4_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[20]),
        .Q(\r4_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[21]),
        .Q(\r4_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[22]),
        .Q(\r4_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[23]),
        .Q(\r4_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[24]),
        .Q(\r4_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[25]),
        .Q(\r4_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[26]),
        .Q(\r4_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[27]),
        .Q(\r4_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[28]),
        .Q(\r4_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[29]),
        .Q(\r4_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[2]),
        .Q(\r4_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[30]),
        .Q(\r4_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[31]),
        .Q(\r4_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[3]),
        .Q(\r4_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[4]),
        .Q(\r4_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[5]),
        .Q(\r4_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[6]),
        .Q(\r4_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[7]),
        .Q(\r4_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[8]),
        .Q(\r4_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r4_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r4),
        .D(WD_IBUF[9]),
        .Q(\r4_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r5[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[2]),
        .I5(A3_IBUF[4]),
        .O(r5));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[0]),
        .Q(\r5_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[10]),
        .Q(\r5_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[11]),
        .Q(\r5_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[12]),
        .Q(\r5_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[13]),
        .Q(\r5_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[14]),
        .Q(\r5_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[15]),
        .Q(\r5_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[16]),
        .Q(\r5_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[17]),
        .Q(\r5_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[18]),
        .Q(\r5_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[19]),
        .Q(\r5_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[1]),
        .Q(\r5_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[20]),
        .Q(\r5_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[21]),
        .Q(\r5_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[22]),
        .Q(\r5_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[23]),
        .Q(\r5_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[24]),
        .Q(\r5_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[25]),
        .Q(\r5_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[26]),
        .Q(\r5_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[27]),
        .Q(\r5_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[28]),
        .Q(\r5_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[29]),
        .Q(\r5_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[2]),
        .Q(\r5_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[30]),
        .Q(\r5_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[31]),
        .Q(\r5_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[3]),
        .Q(\r5_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[4]),
        .Q(\r5_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[5]),
        .Q(\r5_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[6]),
        .Q(\r5_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[7]),
        .Q(\r5_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[8]),
        .Q(\r5_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r5_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r5),
        .D(WD_IBUF[9]),
        .Q(\r5_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r6[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[2]),
        .I5(A3_IBUF[4]),
        .O(r6));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[0]),
        .Q(\r6_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[10]),
        .Q(\r6_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[11]),
        .Q(\r6_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[12]),
        .Q(\r6_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[13]),
        .Q(\r6_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[14]),
        .Q(\r6_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[15]),
        .Q(\r6_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[16]),
        .Q(\r6_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[17]),
        .Q(\r6_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[18]),
        .Q(\r6_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[19]),
        .Q(\r6_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[1]),
        .Q(\r6_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[20]),
        .Q(\r6_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[21]),
        .Q(\r6_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[22]),
        .Q(\r6_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[23]),
        .Q(\r6_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[24]),
        .Q(\r6_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[25]),
        .Q(\r6_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[26]),
        .Q(\r6_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[27]),
        .Q(\r6_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[28]),
        .Q(\r6_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[29]),
        .Q(\r6_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[2]),
        .Q(\r6_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[30]),
        .Q(\r6_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[31]),
        .Q(\r6_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[3]),
        .Q(\r6_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[4]),
        .Q(\r6_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[5]),
        .Q(\r6_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[6]),
        .Q(\r6_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[7]),
        .Q(\r6_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[8]),
        .Q(\r6_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r6_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r6),
        .D(WD_IBUF[9]),
        .Q(\r6_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \r7[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[3]),
        .I2(A3_IBUF[0]),
        .I3(A3_IBUF[1]),
        .I4(A3_IBUF[2]),
        .I5(A3_IBUF[4]),
        .O(r7));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[0]),
        .Q(\r7_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[10]),
        .Q(\r7_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[11]),
        .Q(\r7_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[12]),
        .Q(\r7_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[13]),
        .Q(\r7_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[14]),
        .Q(\r7_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[15]),
        .Q(\r7_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[16]),
        .Q(\r7_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[17]),
        .Q(\r7_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[18]),
        .Q(\r7_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[19]),
        .Q(\r7_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[1]),
        .Q(\r7_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[20]),
        .Q(\r7_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[21]),
        .Q(\r7_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[22]),
        .Q(\r7_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[23]),
        .Q(\r7_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[24]),
        .Q(\r7_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[25]),
        .Q(\r7_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[26]),
        .Q(\r7_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[27]),
        .Q(\r7_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[28]),
        .Q(\r7_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[29]),
        .Q(\r7_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[2]),
        .Q(\r7_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[30]),
        .Q(\r7_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[31]),
        .Q(\r7_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[3]),
        .Q(\r7_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[4]),
        .Q(\r7_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[5]),
        .Q(\r7_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[6]),
        .Q(\r7_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[7]),
        .Q(\r7_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[8]),
        .Q(\r7_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r7_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r7),
        .D(WD_IBUF[9]),
        .Q(\r7_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r8[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[3]),
        .I4(A3_IBUF[0]),
        .I5(A3_IBUF[2]),
        .O(r8));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[0]),
        .Q(\r8_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[10]),
        .Q(\r8_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[11]),
        .Q(\r8_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[12]),
        .Q(\r8_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[13]),
        .Q(\r8_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[14]),
        .Q(\r8_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[15]),
        .Q(\r8_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[16]),
        .Q(\r8_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[17]),
        .Q(\r8_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[18]),
        .Q(\r8_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[19]),
        .Q(\r8_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[1]),
        .Q(\r8_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[20]),
        .Q(\r8_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[21]),
        .Q(\r8_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[22]),
        .Q(\r8_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[23]),
        .Q(\r8_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[24]),
        .Q(\r8_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[25]),
        .Q(\r8_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[26]),
        .Q(\r8_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[27]),
        .Q(\r8_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[28]),
        .Q(\r8_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[29]),
        .Q(\r8_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[2]),
        .Q(\r8_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[30]),
        .Q(\r8_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[31]),
        .Q(\r8_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[3]),
        .Q(\r8_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[4]),
        .Q(\r8_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[5]),
        .Q(\r8_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[6]),
        .Q(\r8_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[7]),
        .Q(\r8_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[8]),
        .Q(\r8_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r8_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r8),
        .D(WD_IBUF[9]),
        .Q(\r8_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \r9[31]_i_1 
       (.I0(WE_IBUF),
        .I1(A3_IBUF[4]),
        .I2(A3_IBUF[1]),
        .I3(A3_IBUF[0]),
        .I4(A3_IBUF[3]),
        .I5(A3_IBUF[2]),
        .O(r9));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[0] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[0]),
        .Q(\r9_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[10] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[10]),
        .Q(\r9_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[11] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[11]),
        .Q(\r9_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[12] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[12]),
        .Q(\r9_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[13] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[13]),
        .Q(\r9_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[14] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[14]),
        .Q(\r9_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[15] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[15]),
        .Q(\r9_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[16] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[16]),
        .Q(\r9_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[17] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[17]),
        .Q(\r9_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[18] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[18]),
        .Q(\r9_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[19] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[19]),
        .Q(\r9_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[1] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[1]),
        .Q(\r9_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[20] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[20]),
        .Q(\r9_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[21] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[21]),
        .Q(\r9_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[22] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[22]),
        .Q(\r9_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[23] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[23]),
        .Q(\r9_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[24] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[24]),
        .Q(\r9_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[25] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[25]),
        .Q(\r9_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[26] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[26]),
        .Q(\r9_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[27] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[27]),
        .Q(\r9_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[28] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[28]),
        .Q(\r9_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[29] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[29]),
        .Q(\r9_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[2] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[2]),
        .Q(\r9_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[30] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[30]),
        .Q(\r9_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[31] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[31]),
        .Q(\r9_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[3] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[3]),
        .Q(\r9_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[4] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[4]),
        .Q(\r9_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[5] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[5]),
        .Q(\r9_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[6] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[6]),
        .Q(\r9_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[7] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[7]),
        .Q(\r9_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[8] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[8]),
        .Q(\r9_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \r9_reg[9] 
       (.C(clk_IBUF_BUFG),
        .CE(r9),
        .D(WD_IBUF[9]),
        .Q(\r9_reg_n_0_[9] ),
        .R(\<const0> ));
endmodule
