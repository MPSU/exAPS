`timescale 1ns / 1ps

module tb_fulladder32();

parameter TIME_OPERATION  = 100;
parameter TEST_VALUES = 3000;

    wire [31:0] A;
    wire [31:0] B;
    wire [31:0] S;
    wire        Cin;
    wire        Cout;

    fulladder32 DUT (
        .a_i(A),
        .b_i(B),
        .sum_o(S),
        .carry_i(Cin),
        .carry_o(Cout)
    );

    integer     i, err_count = 0;
    reg [103:0] running_line;

    assign A = running_line[97:66];
    assign B = running_line[65:34];
    assign Cin = running_line[33];
    assign result_dump = running_line[32:1];
    assign Cout_dump = running_line[0];

    reg [32:0] Sum;

    initial begin
        $display( "Start test: ");
        for ( i = 0; i < TEST_VALUES; i = i + 1 )
            begin
                running_line = line_dump[i*104+:103];
                #TIME_OPERATION;
                Sum = A + B + Cin;
                if( ({Cout, S} !== Sum) ) begin
                    $display("ERROR! %h + %h = ", A, B, "%h", {Cout, S}, " result_dump: %h", Sum);
                    err_count = err_count + 1'b1;
                end
            end
        $display("Number of errors: %d", err_count);
        if( !err_count )  $display("fulladder32 SUCCESS!!!");
        $finish();
    end

reg [104*3000:0] line_dump = {
98'h0f3d496abab877c4293e2ce81,
98'h012e79861ce8db62127d704bb,
98'h073c9ac8392b98870785d53a0,
98'h151a988f751a1eff701a0cd3c,
98'h0e0399e5c7185586f28d2de3b,
98'h01151b896a15da2fe546fbdb3,
98'h0413aab1e75bbc8ceacabd6e5,
98'h183dd299bb8c9b954adbd9cfb,
98'h0f127ec7e4c7015154f29b8bb,
98'h0b3a441534b2463facf660064,
98'h0d21b2758341367dcffb22953,
98'h15320180a41f22b06418ba3cd,
98'h0c0119b8c227f6ab0e54490c4,
98'h0b362c91ac765fd8a38a4418f,
98'h0208bd3cd157fd62edeb231a9,
98'h02192c2cf2530419e4d82ea7f,
98'h0b37875faf36b01d2d1b0c11b,
98'h012b9167172c4e438e9b8ddf3,
98'h0703a12ec7459743c615f7eaa,
98'h05032c85c6528698e3924e1ca,
98'h0e097f6652f8c72ea2d56cc7b,
98'h19a151fd02953fc8e84091a54,
98'h0c269f730d393928270da4718,
98'h013d4f733a9407f56657f626d,
98'h183cf47339ec14680ef455da2,
98'h0c2810bc102a89af148a4236c,
98'h150c0432d807e7184714a69ac,
98'h042df4dd1bd91cf7eb44fad2c,
98'h0d3cb42eb970cf512801c4754,
98'h050bd30bd7bac83fb1ab60dff,
98'h052cc6949984941c4731a6d2e,
98'h0d3c2fac3849b167c7ac56ac3,
98'h0e3707412e2fae7211617844f,
98'h0211a1546362fec18f19ad6cc,
98'h0d2528c10a54423c695d28057,
98'h020365c846eb280d85de5abf6,
98'h0228515210bc0752a23ba3757,
98'h198126fd4263b77d84b916293,
98'h002557e08abe227fa6f9379eb,
98'h1512f01865f37ab1a2b8de981,
98'h0711b10a6371ee7b2ec19ab28,
98'h153a526f349223bb6aa0e7e16,
98'h0c0e0c1b5c37b4eeb2731d8aa,
98'h19b9ba85b3785a1b2a1170428,
98'h021ba010f7505773734c85283,
98'h0a16f511ede53bc20e5afde11,
98'h02392898326ce8918dff0c34f,
98'h181de3f7fbfa4e122d29844a6,
98'h1524930e090f34c355060c828,
98'h1518634cf0dededb678cf1f45,
98'h002e5b7f9c843b70d17dd08a1,
98'h18205e56008bd55f472ca5bc1,
98'h003b99aa373197f2a62b0ced5,
98'h012114890210f34e6ddb4c673,
98'h1983bdfac75eda9360cc81f5e,
98'h180c8e89d91485c9e838a6239,
98'h0c06fe8d4dd3d18a6c484514f,
98'h183a432db4be8662a676b405f,
98'h042a742f94d4c201733e32641,
98'h0c13ec7a67f02c1a263fcd8c4,
98'h0e16e75eedf591112d0106252,
98'h0a258ca38b18ec616f031e1c0,
98'h0f38787fb0d6396be54f9e414,
98'h0b36ae00ad5fd1d67003ac7ae,
98'h022e7c819ccd74ffce259ff5c,
98'h0124033f083f617aa7befc605,
98'h0a30adf1214153594258d92e7,
98'h0d13c2536783c213cadc80529,
98'h0b3d626bbad25c31ed25e119c,
98'h072b759296d80ab27183efa76,
98'h0c0e9a3ddd03b632c780e0114,
98'h150c7282d8ca77d74a44941c2,
98'h0f204d6400afcff40b75ba968,
98'h0d3f5ed7bea6ec7383f407560,
98'h198e688cdce4f8ff92f992d2c,
98'h040fe576dfd7e2e86d9cd8631,
98'h02077a13cec2eacdc8f9f217d,
98'h0b0d9b74db3ece06a43299386,
98'h0f010f06422241c809931a5ee,
98'h0d1715176e24ea0f0448d4339,
98'h0c0ac021d5bee647aeceffc99,
98'h0e042ad348557db3e872699a6,
98'h020ceed2d9ce6594c5966a21d,
98'h02346e4ca8e28b1406f6d519e,
98'h02303236a05b3ae8eac5be582,
98'h0b36cf59ad84f0c248a2db47e,
98'h0f1a741a74ee086d0e2ef006f,
98'h022f70ff1ef8fabeb1021f21d,
98'h0f1ebdfa7d7dc03a284a1aef7,
98'h0b10ae716168637a13271f8d2,
98'h022cb604194fbd594b1e447ad,
98'h042c501618a2c4d686df1cd75,
98'h0a3ccc14b9a0ccc28733c53b2,
98'h0d11f081e3d5792470f76635c,
98'h022616b90c2026608c39da699,
98'h0b1f9179ff23ec2483918f466,
98'h003ae02e35f5560bb290df679,
98'h051960f2f2f15c082d8c0d8e7,
98'h1538e360b1fa148c2e02af3ec,
98'h040dae125b5d0a7071ccbdfb3,
98'h0e0a38edd441109bc7daae20b,
98'h0a3a0e2cb421dd6d8892d2626,
98'h1803f422c7f2a7e3af96fae68,
98'h0e16b1c76d7a7081a7fda701a,
98'h0b3f6ffcbef88ffc2ee448924,
98'h151ce99779da959d728dfffe3,
98'h151b4c27f6a16f6e93bddfcd3,
98'h070ddb815bbf4620b2ef2ee59,
98'h0f211a02021566b468b348688,
98'h0f2e679a9cc603de444da02da,
98'h043cb997b96489350afd1ade3,
98'h011d3d287a6caa158f6850b32,
98'h072266a604e8464b8ee279cf7,
98'h15181f9ef00aae794302ab3c6,
98'h0e30759a20e0c23f9148b3860,
98'h05355ba3aa84d228cbc44df66,
98'h0d09c09153a71f4b0bee8b731,
98'h18066c0bccec42b5882c37f71,
98'h0b15c457ebbdb696293cabb05,
98'h0e08cedbd1aa2b210db4debb8,
98'h0d036d6ac6f7413a27ecbe7f3,
98'h0d3a0a493408b4dbc4feaba94,
98'h001b94f7f71df1407050afc93,
98'h1813e1b8e7da78c76dce618e1,
98'h0b202ddb00737aa12ffb96a01,
98'h0525babf8b71603422e4ea1f1,
98'h012521a20a530c45e425c6bcf,
98'h0d303222a045f5e342de0b7a0,
98'h073fdd8a3fae39078b5d8a017,
98'h0417e0d6efe0270591bb85a46,
98'h011a8f7ff50dd0af4cfe01f71,
98'h013451012882743ccd8a180bc,
98'h0e281320102fa8f60a6db14f7,
98'h0e3022f6a04892994795ef058,
98'h18258eb80b0a5684cb9e2d63f,
98'h041f623c7eda7c9c68cbf94f3,
98'h0706c044cdafd5f410be77b63,
98'h18210a870204f336c52da58e3,
98'h0419fa7373f824cda6897f6f7,
98'h0c10bcbc61786ec9ae0487d04,
98'h0120d1a0018cca8a4b624ae18,
98'h043da3f0bb5f8025e0ab670a9,
98'h198a78d954de51926fe74905a,
98'h180b8a68d72da18c0b9a329af,
98'h0b2cceda19bcb03fabce4afd3,
98'h0f131e9ae63777aea93a5fc67,
98'h01091b11d23ba1daad52a5926,
98'h0a06682a4cd582ad64d12f3b2,
98'h15197a9b72fbef9d25b6fab5f,
98'h0b0e6ced5cc23f1952055a8e2,
98'h0213fd44e7e2a9af09f42b01a,
98'h0a0705e8ce14b6f3ea7da9bcf,
98'h0a00728b40f7502a2606ef373,
98'h052de4511be882ad82bdf0ad6,
98'h0d2de69a9bd1ec17684599bfa,
98'h0f09c68bd3b43a27aa3ff4ac8,
98'h1504cf5149b2186f28af802ce,
98'h023edd2d3dbf55b3a7adb9f02,
98'h0a22e93b85c7fb1acfff8cb83,
98'h00355ffb2a987f11e3fab9159,
98'h001dc496fba82df38ab377c34,
98'h052752ea8e9d52736ef17ca29,
98'h0239024f321397c264f129578,
98'h0d1a7b1ff4d48f796d1326846,
98'h0d0d4102daac3540107bc2a65,
98'h013b83f0370bba34c9ee5d90b,
98'h040cb9fdd95fd215ee11cf893,
98'h19bf53e13e992c26e75b2304f,
98'h02028e3d4501b1dc561620020,
98'h011f91a6ff13954061c110066,
98'h0b19c36ef3bc291cb00cc9b9d,
98'h153759272ebfece22fb57b22e,
98'h1828f0ee91f3265030fdd1825,
98'h003520762a66d2dd0a8705cfb,
98'h0e2f9cca1f20aadf0aa6fcd4c,
98'h1986ccd9cdb260732b5411ea4,
98'h0d2248be84a4342389ce4b534,
98'h0114f7c669e5695404719f388,
98'h07122f38e46e14658abe98469,
98'h0f1263e164ed2ca18ae010e79,
98'h0e2db0559b5fbbdf6cffe420b,
98'h1994a1ff697e75ecaa635b0d4,
98'h18066ee24ce9f1b810c4c5fb0,
98'h001ae625f5df2e36693c18269,
98'h19ba1d5b3421fd0a0d7e85171,
98'h0e180c88f02d5cef137706994,
98'h180afaee55f6bdde2f915a5df,
98'h0004ce8e49a498f80b806e332,
98'h19a500778a1eb62d626a59e19,
98'h19af27cb1e52e9a368f0eda94,
98'h183cbd85394802e04e00845ba,
98'h012beb0417de17b0746130195,
98'h19a4e55289c344cfc64280ad2,
98'h003f872e3f2a6e5088da0a889,
98'h07278bce8f1279c5efda7d5fa,
98'h0702fc6ec5e3ec26058e81652,
98'h0f2012948034c57a2339ba253,
98'h0c3a011a341ae440e3d53603b,
98'h0d02c5f2c5b82a96b0153956c,
98'h0d3f56b5be950f2164aebc226,
98'h0d2f29e59e4a33b452f51975c,
98'h011c4ef6f8a40bb98ade57667,
98'h0f19f719f3f08c5bae7016ac1,
98'h181080c1e102506ad0c2a0dd6,
98'h0b0bc7ecd7828a064e44b44b2,
98'h043ead2c3d678c0488a3947cc,
98'h19a1756b82eca51c90698e4c2,
98'h0d23d47a87b576c9a72386a20,
98'h002b24531676e1f7a53652d11,
98'h002d7b221ace1369c5a88192b,
98'h153702102e3729e126bee3a2f,
98'h19b41ec82814600670db8afc5,
98'h0104b1c04948941150721fb3a,
98'h198edb415d887730429351746,
98'h020e692fdcd09eb16dc5d49c6,
98'h18253f920a6020e887b7c1f85,
98'h1984bddbc94b57da48a1581ea,
98'h011452f0e8acd3a088b4056d8,
98'h150a21f1d44776954a7049a45,
98'h0d2bc9c117902538ea546621c,
98'h042b114e162b63db092efbbe8,
98'h18386a9930efac0286959d4a4,
98'h023fee7e3fcc3395524a05a6e,
98'h0700a33d41494fbed0830884d,
98'h05158fbf6b0f8d9bc2127cbf0,
98'h0b084da250b90a9eac094756c,
98'h15297bfd92c186b8c6f056104,
98'h0e20a4ed01711a42a9fac0ad9,
98'h1536d7d72db769a423e46fcbf,
98'h02396a7432d5a0bc70bb905ed,
98'h0501029842087007cd43c2cc2,
98'h0e183abaf05cb58c61c25ca80,
98'h0738e33db1d56b7c6f9d3c11d,
98'h0d0b1276d603e6a34e4393ae8,
98'h0109e57553c85e8ac8c3be468,
98'h181b038cf61c2963653491000,
98'h050ba69b576505ac138dcb3c1,
98'h00341a11a81d3b9c671c2b11d,
98'h050552bccab35049aa14556b8,
98'h0d27714b0ee1749003ee28c1a,
98'h051fb1977f7cc9bba7023976c,
98'h051c78ae78db05ef71271ed4c,
98'h0d12e397e5c5f24c4f7ddfa77,
98'h073668deacc3acdaccb635790,
98'h0d0cceda599c88336cfe856e5,
98'h19a2e8b285f7d2e3a9aa55c37,
98'h023d3c2cba43c09a47e6aee59,
98'h0536e22f2dde1f0b6f203f31b,
98'h0c24a40b8977709a2cc5404ea,
98'h012e87889d2c76c2056705297,
98'h0232aba4a56f263c0796bf92a,
98'h0b1588246b0b6ee9c9e874782,
98'h0d3151d422ba31792d883dc38,
98'h0a0c7596d8c92cd24bfae0d35,
98'h0229cc2793bd9d3a28b5689a4,
98'h0f1058a5e0bcb73d2579da587,
98'h0f2013db800d1857cbf343f8c,
98'h0e197645f2eab75c03cb4b0cd,
98'h183222dd2447ce9bd0410b687,
98'h0b16449c6caca9cf0f1e7c5e3,
98'h1517e0c96fd231be6df0bb9ad,
98'h18378ffdaf0b7fa7d13a84a1f,
98'h1530bfed2175b268b1d0c3e95,
98'h0232cfefa5aeaf668da99c957,
98'h19bc0a46381f693469f85fd58,
98'h0e0fac265f70b5fcb476dcdea,
98'h1508de80d1a6afa98b601888c,
98'h0c05b187cb5a07cbe9abe38a9,
98'h0a1adcf9f5b4a94225d7ee54f,
98'h051f3727fe7371a42ff3e18f0,
98'h023084be2115bc66f0e4aa330,
98'h0706734c4cd0e9c6e8d190494,
98'h1508408bd0adfb6f84f5d744d,
98'h0e11c069e3a5d0e4896d8efed,
98'h003123cea2797da72c6de4539,
98'h07141225e823a31f08aaa85d7,
98'h022457a488b1a8452bcded513,
98'h07269a548d14190762b57ffa7,
98'h0f1437da68606773050eacd70,
98'h0f109dfbe10fb89dcddd27d35,
98'h198e1fec5c1a574a6c0815a66,
98'h0c227a5004e1d6538d6a1dcdb,
98'h053be80837c8dcd344411428e,
98'h0208d9b6d19b060a6f413136d,
98'h0a02120ac41d2f0764e8f7f05,
98'h0b0d18c4da02fc11c387d0449,
98'h0c27a6808f754fcf29440535a,
98'h0427db3e8f8ade2c46e73d93f,
98'h19a4c1a789abf50384ecae5ab,
98'h0c3ad119b5910489e8d42daac,
98'h0d24d06c09bc616eb072f568e,
98'h0136ab7b2d772acba5b84c76b,
98'h18397d6bb2d32dc86bab7591b,
98'h19a241b784bc110332c32acd0,
98'h022b4df2969501b9e79794aeb,
98'h0c27e6540ff98cb1263013eb2,
98'h0f04eefe49d43cdc67085cc15,
98'h023dec063bd809c6e6364af6b,
98'h1826323b8c5e8fb8ef857d734,
98'h002f5ab21eb87ba42921307d2,
98'h071bbb07f77b84c827b9f5959,
98'h0e39d46db385be1bcfa5cff40,
98'h0e285b6f90a4f973906fe4a25,
98'h1525aa7d0b4e666d47b35538c,
98'h001d21307a728714281d043a9,
98'h0d2d22559a78044a2ea3ea112,
98'h050d12b65a20dbf209e949a7f,
98'h0d37ea9cafccd2d447cb7baa1,
98'h00199c1ef30e04474f412f5c3,
98'h0b1fc026ff94d99b6cc9e8198,
98'h0b04ac374973a33c32ad26709,
98'h182342f8869b7da0651e13dce,
98'h19a5817c8b181beae7afb0264,
98'h181bfb4877f28255292f6759e,
98'h0f0d271b5a5faa5a74039f676,
98'h0b3c8e79b9337a9aaa5b345d7,
98'h0017a1f16f566c85711c02451,
98'h198c2422d870a9c12bdb839db,
98'h1996cd8a6dbc5b542c7f33790,
98'h0a03fb0747f6548ab1d4ca37a,
98'h19b3e92427cc33a0447e93e48,
98'h05242e1d886d8227106007311,
98'h0c14d4abe9a64f3183646c112,
98'h0c04a989c9612d380d6ec8f75,
98'h0001fdbe43f86dc2255975b07,
98'h0b174fa16e96e4cee0fe9ae02,
98'h0c39fca833eb6dfb0e6b8d1c1,
98'h0d004de9409bdd6bf0095aa8c,
98'h050fe166dfcff674c3670ad55,
98'h1519a216735772006937f5f6e,
98'h0c2130a702730eb8321c4505b,
98'h0a26cf0d0da414ec83a50fd7d,
98'h072090c60133a83e25f2b8fe6,
98'h0a2dc1e31b9fb10362150e411,
98'h0a2226d08462177089735cb9a,
98'h0a19e6ddf3d47a83e3a10f904,
98'h1506a3844d627ca80f7b98587,
98'h0c3e6e71bccb3020489a480b1,
98'h1812004d643b1d2d324267a47,
98'h003cc2433987cbf8cf13475ea,
98'h042aec4915e7ac390e71238ef,
98'h07042a284861a49e8684a6208,
98'h072fe9449ffa83f5a3d973b1b,
98'h020fa125df57fe1369ca9b4e9,
98'h0d3f18bcbe04ce7ac859e7ce5,
98'h0b36da6fadb40ac6b2d0f9cdd,
98'h013db8debb6e9ed18e3ab94d9,
98'h0517766ceef95c9b2f2b15ec0,
98'h071c51877897f9f36d0434c20,
98'h010b67b056d5c5e0efed12deb,
98'h0c049143c90bcfc945f84b645,
98'h181188006331aa59254418434,
98'h0e0dda50dbbde42c2ed0cc966,
98'h073d5d513ab1c034aa72ef9f4,
98'h0d057f9b4afca7e4b07bc7617,
98'h0b330ec8a62b4114860089e00,
98'h0a07b1c04f7001ac2c5793f74,
98'h182489bb093b8b0a265decdb2,
98'h0a161c0d6c2e072c085805315,
98'h1834d6ada9a431960d9108ce5,
98'h0c09317f525ea5fcf0764210e,
98'h00169e55ed3c7ea9a799f5df1,
98'h012929c212573ca76b54c73fe,
98'h0b2ade9795b963a524e0199a6,
98'h022bae34974723a4c839108f3,
98'h0d14cf8969bcda5aa65cb4765,
98'h040336e2467e265dadb46a790,
98'h0d27f86e8fcdb60a42a057500,
98'h181d1788fa05ec2c473d6b9e3,
98'h198574bd4ac8e465d488c0ed4,
98'h071b3c94f677515829139648c,
98'h0c2d691a1acd1e8d4f64a37b4,
98'h02069823cd24b01b89bea1e9d,
98'h0739a85a33520a1263cad20fd,
98'h04273f020e62199e8ea2ec9b2,
98'h0a2688820d0bc9f5c4a256282,
98'h051f35ad7e647efa85cc949df,
98'h153ee7c7bdebffa810e0ed29f,
98'h0014ed5269e0ca3894cab9dbe,
98'h0f30618f20c13c0bca7d6de2b,
98'h19aa70cd94c3e751cbfc6766b,
98'h013cb36e3965e0708b9b9607d,
98'h182e41ac9c8cbd2e4ea8a4f7a,
98'h0f2d52291a9f6f97ed2ebfb6b,
98'h0e22e52c85c116a84a7330704,
98'h0b1e2eb57c7f4eb224f8fef53,
98'h152a213a14667b8791e75f59e,
98'h0424ab378945f6614a6427306,
98'h0e10e972e1d7f986e35aa8663,
98'h0107c0054fb993b5abfa38be7,
98'h0128fc2291c1dd4d443054eec,
98'h0c2e50a29c911930e4bab65bf,
98'h010d2f475a7c5b74aa2fda74e,
98'h1998b0c5f144bfc346e262af0,
98'h021d6d8dfaee298612b75c224,
98'h182a59529484f7ce4f42e5c4f,
98'h19af63529ed006faeb2bd4483,
98'h0c38cd5f3188ca224e1fda936,
98'h0520dba3819a363aef7065e05,
98'h0104af2f4954a900e1aec477a,
98'h0128cd3c9194e5a06296560c1,
98'h0a320539240ab11b44af6cb74,
98'h0034178c283488732b8f2d951,
98'h0a04af20c9455a91ca1a27ffd,
98'h0b0aefadd5db1fede4d2826ca,
98'h0e160abbec2d99f5883983e6f,
98'h002bfd6f17c77437ce90e92c5,
98'h0528c90f11ad714805fcdc69b,
98'h0c3a284db46b3d6a85b58e95c,
98'h0c2ff34f9fcff0fa5029596e0,
98'h050a147554113c8feafff9127,
98'h0d0e1fe25c0fa8ec4646d4415,
98'h150c4fc3d8ac449f8a477233a,
98'h0d01d75bc38489704b6e2518d,
98'h19812ec642583383642198330,
98'h152429818852344666f658927,
98'h051359b96685db14475d97720,
98'h0b0e72495ce7bd9f8ae64d336,
98'h152609898c3ada1aa9fd8bfa3,
98'h182c4ed61891dd1de85838e91,
98'h1813f4d567fe6550ac2f8afd0,
98'h042ec27e9d908ed1700496898,
98'h150bece857fc005e286fd4540,
98'h01058bc7cb11243b6b41fb51a,
98'h0c282abf905526dce305ac00d,
98'h1833a965275dc54ce71f54672,
98'h000d4c095a8ae5554fe45bac8,
98'h0a040f3dc8036166c6a60c57a,
98'h180e00215c186240e481dc292,
98'h02138b64e71f1059ed0998989,
98'h00006514c0c75707ca4ca6efb,
98'h1514db2069b3e367a031ef072,
98'h182214a1043779042fb22fa20,
98'h0f23efe487da2640e71663695,
98'h0717e1336fc1d27e45bf85896,
98'h152d64579ac910064db66cec6,
98'h010642e84c910bafebfd9d177,
98'h021f214dfe6be4490365d3a61,
98'h012f748c9ef7a3c0b022c165b,
98'h050732cc4e63840a8809c6135,
98'h0134409da8bd19caa4daadb5b,
98'h0035cd072b856ebbca7c569a1,
98'h15047e48c8cb05d6caeecef0b,
98'h19a781648f19333ce773e107e,
98'h073c3e6a385321ddea302d286,
98'h022ca379994550dfcfe3d8120,
98'h199aa88ff57742c8a6dc7d165,
98'h1532de0aa58c8864d3c47ad62,
98'h0a2f87f51f2c41700eafd99bd,
98'h1985f80ccbec9cfd0a56f2594,
98'h150c88895900d39e495ca5427,
98'h150cc9a5599f854aeb835709e,
98'h183723e72e61550a8bab13bc1,
98'h15376128aef00c5d31a61e3c6,
98'h0d083e5d5061805f1109db617,
98'h0d03581c4682e2b5c75a6faf1,
98'h151673e86cc51834c4e18eb48,
98'h012b583516a51f461076e3074,
98'h0e3815343030801425f41ddec,
98'h1506d0584da1306f0f9a25521,
98'h1519d49f739a4576e8aa0031d,
98'h198ed99add8b3d01522d06859,
98'h0a1723366e4698c54dc685a70,
98'h182d4c411aa5f53e0e176efee,
98'h15313db5a245b6584cb4d05fc,
98'h072b04c09630d3d62dddbd037,
98'h0731e98aa3de3f79e756f625b,
98'h150258bec4a0ceea8ac40a412,
98'h0136e1d2adfc8361a668c9ea5,
98'h050abc0fd574790cabccd94d1,
98'h0a12f45a65efb839869fcd472,
98'h0b2295b88504923d4c00ab24f,
98'h0021ce9e03ae241a8409c9fd7,
98'h182c44ef18a208ed00f3fcae2,
98'h011b7acc76c9360dcc3393770,
98'h19a3561786826afd4df92c368,
98'h0a248cc0892a8f0b880970453,
98'h183ee7c7bdebc6bf04d3c6f30,
98'h0507ff08cfe2fafd958aaba1a,
98'h18063fc3cc40fbf3453abe819,
98'h0237bfe1af4459bc4911ceedc,
98'h0f2c9000993f7ccb2c5f06677,
98'h0120ee3801ef78110a1b0332f,
98'h0e38eba3b1ef7ee700c419924,
98'h0410c6a9e1aed8b4900a1aa2a,
98'h0a2f6c029ef79c58a96fe7d79,
98'h00174082eea76d500a49c216d,
98'h0e2085a10134e4a0abafab74b,
98'h07045ac048983f7ce3d55a907,
98'h00338d3527285daf83e7268f5,
98'h0b0d190fda1209c369d6fab92,
98'h0a316ca322faf4e7a947c8b4d,
98'h071530cdea7fc09cab4b1862b,
98'h0e0488004908e018cc653c5aa,
98'h0d0a660754c90b7245c35a064,
98'h0412d291e5956e84e874dc5e6,
98'h0c2e98799d07ad9c4a6a1045b,
98'h0a0713ccce3849dbaa4d91857,
98'h041d80927b38df64a60fd76a2,
98'h070e5c555c85273f4fd597fdc,
98'h040b1c6cd6039703c8e4e0e52,
98'h0b3eab013d5ee8406683acdc2,
98'h0227ccd70f9cc1a2f22764d06,
98'h040bc1d5d7972bdfe471239e8,
98'h0e07224e4e426c5ac6e8bb6d7,
98'h041f2b077e6b4f8e871263aa4,
98'h0b1659ff6cb6dd34b0a29ea57,
98'h18186dfaf0dfe02e6df34dcd0,
98'h0f1f8ac6ff149c29f23e138a5,
98'h0c2a744514eb7b0e938d09bc3,
98'h0a0682324d046c22c8457bd4e,
98'h003b1eac36121ef1e5c2bb954,
98'h001c517e788e33f84d934f678,
98'h0f1a0a247401ed08ce2aa15da,
98'h02168a97ed2dd77410c6fdcb4,
98'h0f1384d2e73259f3abd11882f,
98'h19a72d1b8e45004ecd9177b1a,
98'h0514b30c6976cec429fb0b5a9,
98'h0422435784b2d7312ba2e0742,
98'h0b05e4564be5b9fb023546a23,
98'h070e2f48dc4aacb4c5bae7945,
98'h0a301864a025108908d636ff6,
98'h042ba79b175292626a954a3b6,
98'h0c32b41e255d3ed066df8e7f6,
98'h0f3264ac24e2e3b28c63fcbba,
98'h073e66963cc389a0cd055217a,
98'h022f7d889eefbf0f11007c0db,
98'h073a3e12b45cdf3b6847cf25e,
98'h0f2274ee04f56ed02ee5c7538,
98'h0527ed080fca18514505f8ef9,
98'h0c25f6490bf0c23fa53c81565,
98'h070c3f1c585ea903e605ae223,
98'h052142b702bc5695a7daba081,
98'h1990be236172c1e3a1f766533,
98'h19af4e049e9bcffbeec0e001c,
98'h0a0387224711e0f26e12c7802,
98'h0d188baef12e028a84455a053,
98'h180a4f4ed496d2a06f91a38e5,
98'h152c6be298ef0b4b8b28487bd,
98'h050d990d5b3622ceab86ddcb8,
98'h0b37887d2f2359378810eef70,
98'h071118f36227fdce0e96b86d2,
98'h0d03820b4734a637aa4e45b05,
98'h0a1e4ac57c928160e50e0a10c,
98'h0b3d8cca3b39e02431ac33099,
98'h021636786c457db6519ddb3b9,
98'h0a10ada6e15301c76b96ed0ba,
98'h0d2f65319ec8a6704ad8ebdb9,
98'h0130a73e2171dbd8aafe02e87,
98'h021506466a2d339f88a8a0c5b,
98'h070296dd4518ce026b108e797,
98'h180c443ad883f2c5c306d937f,
98'h07004180c0886fdccc240dc02,
98'h0b34c9c4a988c7d341e22c576,
98'h0a2310d6060529f14d2f6465f,
98'h012976c892c49e28c40a0eb1d,
98'h0d13c03a678dbeb8c4fb853c5,
98'h0c36455c2c96c9986d285fbcc,
98'h010bb9ba574bc39c4e3343bd2,
98'h00085ec3d086d761c615df55a,
98'h19852312ca7709f4a423cd896,
98'h0b2d60741aefcf3688ff0b41e,
98'h02069ab0cd14f80ae9874beaa,
98'h0126d1130d85e438c3c6e4aef,
98'h0a07a4b14f6cd21783ab2d52f,
98'h0d06c5754da795f7865d1db23,
98'h0b1ac7e1f5b9f344a6ab96db3,
98'h003ab59f355b4174f0352ec9a,
98'h013a5abf3494f6ab6d657dc50,
98'h0f1981c6f30a2221cd73d45aa,
98'h0a050075ca3cd052b088e8fa2,
98'h0c39a7503379c2df251074322,
98'h0126d5e38d98d635efecda8bd,
98'h0e04a5d14974defda3afeb066,
98'h001c4e94f8bcb93ca5de6133c,
98'h19ac940d9904b33f4e3641f46,
98'h0f2bc1c697a76e408cac51d33,
98'h1818e4fc71cbbed3c9b4cc01c,
98'h0b22a7660566070a127928f40,
98'h0c0f5cc05e82f45cc4222b9c0,
98'h0b138510e7337b52aaa494474,
98'h0f0e35afdc4a5aeb4c91c018e,
98'h0b018b12c31e61c3ead62426c,
98'h003c754fb8ee1f000387fb35b,
98'h0b16e1696ded98f50e4aa513e,
98'h0c057154caf1138cae411e979,
98'h0f32a4c1a56ce07085bda1386,
98'h012484a3891da2f16d27e14c8,
98'h020b9378d73a61aea29089e54,
98'h0515f451ebce2fffc6517d49e,
98'h05146a9b68de29196c3909146,
98'h199204a4640de6f84b7ca4ed3,
98'h053ef2e6bde48f088f67fae72,
98'h01273e100e62fe8c90c8e07bc,
98'h072abdc7956490c583e28f272,
98'h0738e239b1c368dd4723d3a34,
98'h0b3c925bb90b1989ce3f12c5b,
98'h0e1690f6ed24f47b1111eaf95,
98'h070b8a6f57343b7e2ecee15c7,
98'h0c121d4c6409dd67c78ff17b6,
98'h0200df7f418b58bb4c06fead0,
98'h0128926e111ace1360e30e0ea,
98'h0a3767b92edb3c4a6490d8206,
98'h050368c346cf505fce44a900e,
98'h0717c2f9efa7232382f4ae48c,
98'h1506eadecdd5ae9d6dafb9875,
98'h0c1e37ce7c55b531e8b7265f1,
98'h0c12ca86e59b448df21cfb401,
98'h0b2740730ea6ee4c8c6b83c53,
98'h0109e5afd3c6406146738bafe,
98'h000fc7d5df9df73d653409844,
98'h04263b7f0c61d3b907eb6fc4d,
98'h0a2616928c37eebca42203ce0,
98'h0b0e1149dc2dd4a685978153d,
98'h0b186ff7f0f8a274a9cef97c1,
98'h050f47945eb2ceaaaf04449b2,
98'h0b3e5f01bc8637fd48f0858fc,
98'h0015df146bab83b611f125bfb,
98'h0b09b35cd37cc5dfaaf058b29,
98'h0b22adae0544dd29c7a19e4f2,
98'h0f1c2e677852dc956419e2b5f,
98'h0b374377aea54cd711dbc2bf3,
98'h002ee02c9dd7ff866e772413a,
98'h151bffb577dc9dfee781b7ecc,
98'h0028346b10460e0cd33e276d1,
98'h199555dbea8d3652441b909df,
98'h0a2daf8f1b4e9c70d108a30b8,
98'h070d4290da8fc6f1c95f12fff,
98'h0b2e5bb61cbd3cec28674260a,
98'h1825f0a88bc26d6ec9fae6289,
98'h0a12e5ace5f7b8a728fa1785d,
98'h011a8e28f52444ca0c02a7950,
98'h053069efa0d538bb6d8fb4bcb,
98'h0e035146468e6674c98168aac,
98'h198af1acd5f55f3125246deec,
98'h1801ad65c34b5b504be014378,
98'h00249fc00930500226d3422d8,
98'h0b09b81cd37dfcad22553bf09,
98'h04068db74d28aa1687a1ed328,
98'h0a2dbe2f9b78c54c244bcdf37,
98'h042058cf00b87048a969a0def,
98'h01010893c216925ee1363245f,
98'h020b5ef4d6a1e26000c5e6bcb,
98'h0716d16e6d95d485e62b50553,
98'h0e2eabc51d5d46176d2b297d1,
98'h0c126913e4e730d20ae2fc772,
98'h0f30958d210ca015cc3e66797,
98'h0f2d8b091b1091c56c0f4d68b,
98'h05130a49e60e5cf54a8f8733a,
98'h0209e30453f5a84faac859cfc,
98'h18078ca84f17ea3ee57fe2d50,
98'h1512c1e96586dcd2c9c7ddb9d,
98'h0037e1052ff13f6b2ea667af0,
98'h0d2402cd8807b01ecc0a481c1,
98'h19b06a6e20da56e3654aecbb1,
98'h021b1ff5f60d8c754ea2b0546,
98'h0109379f52539700ee0a2b1ac,
98'h0d2777d78ec80687c4d733a81,
98'h051ac006f5b22b0ba6fbdf97d,
98'h071ec2177d938e766eb33ac4a,
98'h0d3b50c036994c3e712c94237,
98'h070ab48a554790d250f5273fa,
98'h05322999a4617ac0071491572,
98'h0e14d835e9a1079c8a64e9166,
98'h0f3d4a103aa6a6ab0ded77f49,
98'h0c258e4e0b1a7b46f278fc2ec,
98'h0036ee4fade6490805d002654,
98'h073b4538b6b273b0ab874dd5e,
98'h0017bc366f466cd04f7b6e3a5,
98'h002edd8a1d91592cebd78a41a,
98'h0102a050c54ea7ebc7700dadc,
98'h198a3f08546fc57a8194520f2,
98'h15375adbae8c0434cb7e8120b,
98'h05061da7cc0e44cc50f0d7c41,
98'h0f38bcc43148d8734445189d0,
98'h0a33ee8ca7ff86c23020654dd,
98'h052394a7873191612c8cdd53b,
98'h15090d0d5235ff6da31549823,
98'h0d234bd286af6aa689cfc31ec,
98'h02300fae2035f84fa4f4ad9e4,
98'h01213342027217dd289981ff7,
98'h0f354d23aabd115920e4d2c7d,
98'h19bb80a3b7115d8dee7c979f3,
98'h0c139154672031eb1433378c6,
98'h0a00fb53c1df9a316cccf0cfd,
98'h0a1602536c10e9d662f825615,
98'h041e595f7cb63f302d89bb0a7,
98'h0c343566a86b425c10352623e,
98'h151a4c83f4b539e4ad27ddf0a,
98'h19bd74033adcff2d7273e19a2,
98'h0f2d3f2d9a5e4c96f5269ccc2,
98'h0c1830ce70674f6a8a62e2f12,
98'h0e31c17aa3a557800f1fe00e3,
98'h150aac9c556beea58c75c63ea,
98'h0a1aa637757e91c92a9da6d07,
98'h0d31cb72a3a6b5df0fe64e002,
98'h020bcfe057a3b28b0c3620546,
98'h013b1985b6249c88066be09ad,
98'h0222ada3057909cf2dd7ed836,
98'h0f27003b0e39298121e6eddc9,
98'h152b685c96eb898e07580a6f1,
98'h0a082b285063541c0b05bc7aa,
98'h0e2fbf9a1f50beb1669adfd11,
98'h15251d110a02d5194b601f92e,
98'h0c3c9697b901ba10c7c9fc8a9,
98'h0510f4eb61eee7a9914f942a1,
98'h0a2b31439659e976e9bff7253,
98'h0b0062dbc0ef7a6f082146aea,
98'h0c2b21399672e09b22fbf752b,
98'h0e0fcd375f89d079c8a780753,
98'h0a39e2c7b3e612278b66676c4,
98'h0b1fa582ff41924a4f87fd3bc,
98'h072529ea8a4d78b552984df34,
98'h0b1bed73f7df4ed2e45ca8a7f,
98'h0124df4e89ac2fcc90becf11b,
98'h0033ebeea7fd6c73a2b443c6c,
98'h0a09cd51d397fce76a0c56189,
98'h0c3712092e0c89fdc768728e5,
98'h012dfd009becc86d8e90e701b,
98'h013c1007b8304fb2a746b15b8,
98'h0503c318478306b8ce5b17ee9,
98'h0b271a5f0e05b042c321b2744,
98'h00107d0560d21112664b32a87,
98'h0f145eb5689399cf6838a385f,
98'h198ffde55fd76eb26de9fe213,
98'h051ba8de775716e96e59db25f,
98'h072dab849b4c0dc24f1caff1f,
98'h0f1237df644bdf91c89e6e51b,
98'h0e304b60a0a06c5b0cd785dc4,
98'h199fc2edff825a39cbb42deee,
98'h05257fa68ae8b18616488749e,
98'h0c2bae6e17440cc1c4038c4b2,
98'h0109f43353d1b63c68dbeecbf,
98'h071770f66ef77d7ba536ea9bf,
98'h0f1b3b937667fe660d83bb9c8,
98'h0d2b284a166484279160ce7e5,
98'h0b305c0420a9a1dc88e3eb1c6,
98'h00095e5f52aa0af78af67f782,
98'h02260c728c0c2569c4acda55b,
98'h002efe5a1de63f8b838c8c771,
98'h0c1ba17c774f43c547854f796,
98'h0f34799128c233f550dab9506,
98'h0c2daa6d1b65a6988dfdab619,
98'h04351c87aa01efb549e4d4416,
98'h150b3e42d66c8f7d0b8dc30f3,
98'h013193f3a329f0bc0addf36ff,
98'h0c32f8aa25db70fbe916e12be,
98'h0a32a1b9a57b1c6c2c839a698,
98'h0c14a7006944778d4beb6f897,
98'h052101ee823620952d5647a36,
98'h1984a551c96f029a81d5c8a0f,
98'h01377fd82ec7447948bce9fb1,
98'h0c1deb5c7bc50d7ccbffb1145,
98'h0c243aeb086ba9c811f8be364,
98'h0d1fc98cffbc887d2523f92cc,
98'h0d1e1bcbfc10fda3f33714828,
98'h150455ff4895a1d4724bc65bf,
98'h0b23794f86e0999c87667df4f,
98'h153c8981b936feab248104bb0,
98'h0106ed7c4dd714b4739ce20b3,
98'h19af0c909e20e41b03b7808c3,
98'h011f5a85feb9445b2df3fc2ae,
98'h0c06b459cd60502d0ff627b84,
98'h15201fd10027ad728659c121b,
98'h198dafb95b5b02da6551f350e,
98'h0e0e7ef3dcc1654b4d3a2ca4f,
98'h0102643cc4fd770b2ab3f90fc,
98'h19b930b2b27762a6217ff6d20,
98'h0c02fb20c5c3cb98d30c24d63,
98'h0e072a02ce613eb50471b1ae6,
98'h0d1c9e5279069c4cc71a1a2df,
98'h02229109051466187188cea7c,
98'h073b656e36e4cadf01cdbdc86,
98'h0f34e21aa9eeb9e08f880c134,
98'h0227f2c20fd337f9ee48e6fec,
98'h0c1944bcf2b5a08fa47ecaaf0,
98'h0b2fc04b1f8b6c354fb3b9532,
98'h0e1a10a3741a8715eaaecb201,
98'h05051cb5ca02311ad08d25ee5,
98'h0f3e82b4bd25d1d483c1d3742,
98'h0513d85ee7bf1a23331915224,
98'h181da204fb793d9d2b34bca08,
98'h0037a2532f5dfdb7f4e5b7e88,
98'h181b54d9768ab0afcbe56802c,
98'h0a311550a2335e30b3a981624,
98'h1524a5a689687bbd8b191ce05,
98'h002674c38cfcc2d827a348590,
98'h19b03812a0480ae84348cde6f,
98'h0b2d19c99a3600e62e7e10beb,
98'h0d37edf1afd006c06958c6abf,
98'h0708902f511c74846f41fd2c8,
98'h1990bc48e17ee546a609412cf,
98'h013c637138d929cb6ec3e863e,
98'h0d35b04d2b7eeaecae85634f2,
98'h003d9bbd3b3af5c42e2d26ce7,
98'h0a0b2463d6689b930ede24605,
98'h0400eaefc1d97f68681ceffdb,
98'h000f2521de649b8a81769a961,
98'h04128995e52a38a0079cf02b1,
98'h021c064bf80e00954a4f308d7,
98'h0f14c3ece9804744ce8a81b84,
98'h0d1227d6e46612e28e2542cc6,
98'h023236e124605e1f8c5e0eae5,
98'h0c2deae81bda7e14e9a4a5402,
98'h1500bd10c14185e94a021a3f4,
98'h0b3ed6d4bd8ef23c459090be8,
98'h0d020bc7c403d64ad23372443,
98'h0d24ee2109cb34da44417884a,
98'h041f00037e161edd65bc08bed,
98'h18293383125ea1dff08d47b83,
98'h19aa9b7095338029aaa1f558c,
98'h0e365edf2cba1cad2bb786e69,
98'h0029b16c9351f4a96ebc1ee31,
98'h19a6c24a8db17114a4dee9858,
98'h020c4404d88ac9c4c9d60cd7d,
98'h0b0c5f0a5885245646a5c3726,
98'h013590f52b3608d528e460d82,
98'h05082a92d045b6234b1ae6729,
98'h021fceab7fa1d0230553782d8,
98'h02358389ab11519d707067b39,
98'h00189943f13e9be82b51b549c,
98'h041ed6c3fd9cee546c55cd4b0,
98'h01030f8c46097f4d506ef1461,
98'h0720744580e9e14901c323b66,
98'h073ca001b96d4d6b82029563a,
98'h198e94455d38ddee302a7b5b4,
98'h043185d02303b24b4db1dc8ce,
98'h07238c26873b6723a9cd4e06d,
98'h041df5d67bcf3be64397bcd29,
98'h182b337f9674b03a2ffb4c6f2,
98'h0f28fb9f11f753252ba7f8ee7,
98'h0410791460eaedf3884813b11,
98'h0c3606692c3f24e1293ed9c1f,
98'h002227da847a17802e1d4ad29,
98'h0f3a2620b4607ae281270fd6b,
98'h0013dbf6e789178150e6a840c,
98'h0f11f86363e384e309e73cde0,
98'h053027be20526d07ecbd5f519,
98'h0c05457d4abc918c2960a5318,
98'h0f20e8b601e13c9485b075c26,
98'h00154d6beaa8b77584408952a,
98'h0422cc930593d1196aaf81385,
98'h0722c4dc05b26e29226da76b2,
98'h0129063a12248cf583354cc15,
98'h1528822b1137171f24d364cbe,
98'h002632c00c6a4afc0997e6529,
98'h0237da65afb676c1a3241f6f0,
98'h0d1f6e6afef12f6cac7b9449d,
98'h0d13ae4967651d6913042775e,
98'h0d1e99aefd3ce8f92d1e32ec9,
98'h0d3727422e6ac05e1296e0aa0,
98'h0008ce3051b561c1aee879e80,
98'h0a05246e4a6582da046f8bfc8,
98'h0f0e03c55c2ee057851aa9d21,
98'h000d5799dabb2f06aacf39073,
98'h1816e572edee98bc06b221a82,
98'h0d041241c8315efbb1815f8bb,
98'h0205d66ccbbcad5fa54d5c4f6,
98'h1839c293b3b595c2a370a0f32,
98'h15102719e044a02452fbd6159,
98'h150f206c5e6e48540d5531cf8,
98'h07247a0d08f53359acdf5a301,
98'h0a130a58e61dd69a64066b59b,
98'h0703590d4680bac24c0c383cd,
98'h152712958e10746d636104f3e,
98'h0a1efa0e7dcedc8dc8cde1c0c,
98'h0c37bc102f7e0295b1fb75a70,
98'h01073435ce60c25d8eed6fa97,
98'h150567654af8d7cd23d9fda4d,
98'h0216a4d86d58ba4367ff8fcca,
98'h042aefe215f279bd2bdbd7c6f,
98'h0a06047acc0647bf46875a67d,
98'h183ef8843dcf45fdc583130e8,
98'h0c3aabd2b547a4c2d5838fa07,
98'h001ce8f779f20b18306094255,
98'h199548c4ea81b2ae4e83bd03e,
98'h0b129a99e5189185f105bedcc,
98'h0a35c3662b9f5b53ec0acb07f,
98'h0b1fb5777f5214aeed7547ae8,
98'h0e1952fbf2b961f3329c72899,
98'h0423bd4d8748abed5034ad3bc,
98'h1827c2fa0fb7a43ea2db1a4eb,
98'h0a07ce89cf86a38949f7d9ce3,
98'h0134e80729eccb5606639c84c,
98'h0c210b488210c5bceac86cd74,
98'h0e2b44f7169d6ccb638c74416,
98'h0038b857315e93afe9322c70a,
98'h0704dfcf49939b9eec65d301c,
98'h0c170a326e296e7b84261edb9,
98'h022746c48e8fe9414e901e2b7,
98'h0a1da2077b7bb029a42dcc017,
98'h0727c53c0f98d694f166548c4,
98'h022ebab29d58b4b2e5b026f44,
98'h012cc8cb1999b4e9e7e1dbd96,
98'h0c0e05c1dc06d2ff46b19f6d4,
98'h0211763662f1f700aa0536304,
98'h0e183871f07445e92940db4dc,
98'h01206e7200c5f20b4fa31f96c,
98'h0a1e48af7ca005388079981f5,
98'h0f2ac3a495920eaa71af9379f,
98'h0d215a17829f8ea7e92f3493c,
98'h0d301e22203169eea3f03a2fe,
98'h0e1c5af7f88a9ede4b5862043,
98'h153d116fba38e659b1a9be758,
98'h0738514c3085da75d3dd7df25,
98'h1994a142e977acdc2def8af07,
98'h0f3857c2b09566f770c31387c,
98'h0429f67f93de1dd76ff36fae8,
98'h0c1a4ab7f49073dbe6020515c,
98'h0c1f443c7ebc321b302aafa4f,
98'h0d192538f27eb38bb2b6dd95e,
98'h042edcbc1db84be9afe5f6312,
98'h19ae0e019c18c4616879ca297,
98'h1813767666cf77f44d71b498c,
98'h071d14817a1489a46fb8bb9aa,
98'h1534a10da9601e5a904c67897,
98'h180a9dd2d516748eefa52fda0,
98'h000c6a58d8f023aeab4844987,
98'h198681c44d10bd48e63f2381e,
98'h012b335c164f79f149a5cfc35,
98'h1829d7d293898bebc5deab535,
98'h072eb54c9d6821930aecd8ef9,
98'h0a14742a68f11180a925b5b7e,
98'h0e31368f227c9a752cc1616ac,
98'h010714a8ce2091008c2b74411,
98'h0425efb88bc5c4e943c9e96a5,
98'h04073ddb4e4b585443faed287,
98'h0b07a08ecf5132af6494a58be,
98'h0529c7fe139aa955669634cf9,
98'h0c2e55061cb0e7f8a6311c54e,
98'h18111bfee21d92cbea37cf3fb,
98'h19915a4362bd8c66ae8babb2b,
98'h0d1c207a7865b9718f13b9aa8,
98'h152a639b94dc0c0a7160767af,
98'h0232d6bd259a10ef6a819be98,
98'h011edf94fda7a86409f339eb2,
98'h040da7c4db7884ddafb1a1fe3,
98'h07047ce248d17965e7e18b28a,
98'h0e04613e48ef91c603f57d921,
98'h0a05df6acbb65e6fa5bcfcc11,
98'h0a21e28603e8ce21856f0f76a,
98'h0b1c8541f91c5f52e382ac29e,
98'h0e2979a992cd6358d10e39253,
98'h0a04dbad49b87d50a83db7409,
98'h152af06615fd76c524ef563f8,
98'h01018421c30df419caca19cad,
98'h0a32492824a382af0103de0ee,
98'h0232c944a5a7eacf0bb572f5c,
98'h0c102c0d607c9f50a9f6ad04e,
98'h043743eaae9e95026b2332d78,
98'h182803e1901ebbd1ecb5763b4,
98'h0b3ab0193548c3b3ca11afece,
98'h1820cb2281b5c74bb020dcf33,
98'h0e07f2044feae6548675a49b9,
98'h0a0588fdcb20c9c7877cb6163,
98'h0f234b1186a47bc5854994b15,
98'h02127e4f64c7ed3ec571f1b5c,
98'h0a21bed6834cf358c9b69ae38,
98'h011c02a4f8347699a35bac8bd,
98'h0b22a8178560fdcd8e541e4fa,
98'h182c113a1823aeb10420e9794,
98'h07007dc9c0d14e566c13effac,
98'h002385fe073dbb4f21f473081,
98'h0c3dc8123bb3cb93a1d850535,
98'h041c0a8c7809682bd1fc64e97,
98'h0c234545868830964f095cae0,
98'h0737b3322f65dff004aadd76f,
98'h15343ee928711ddeada764c88,
98'h053b4bed36835535cf695731f,
98'h010e0eb25c329a5f2eefa848b,
98'h0d00556940839b8547502a446,
98'h0c37d3852fb704782360fc3ba,
98'h19bbb204375bb057eefbb5ff5,
98'h01175677ee8b72fa5445d8970,
98'h180602cb4c3f34162be8b25c8,
98'h04301fce2034862729114db86,
98'h1502b47ac54ed3194919297d5,
98'h0e01bbfdc36ca8af069461e50,
98'h0a32bc7fa5729eaaa45b992b3,
98'h070a30abd44cc0b3cbe956ca9,
98'h023005f7a0395602a6d5bc57e,
98'h0c21a1ac835050c5e89a56fe9,
98'h0a3e8eaf3d059f4ac3dc7c9ca,
98'h04142605e85608e671d10b7e7,
98'h0c1034236042309bcb1a8bbb1,
98'h0d0eccec5dadc7860b14992fc,
98'h0e0830815045e8fecaaf251c9,
98'h0f24d2c489b50a86279386600,
98'h0f3b47a5b680d96cc6367752b,
98'h0d2206248432d038316f08449,
98'h0f19a41df37b3dcea45535973,
98'h180f5cd0de93e85c70a5387b2,
98'h0e1f6426fedf65fd6da8d14b5,
98'h0d3eb8bdbd58b524733fb2891,
98'h0c18d6ad71b78ec232a5db788,
98'h0d22dd1085b55c302f74195be,
98'h19b7684eaef8aad5a4b60e503,
98'h0128931f91156791f22c04c91,
98'h0524405788a31be1048f7eac6,
98'h1535ff6e2be3d6c98371d70e2,
98'h0a2d8dc51b325b7db046758de,
98'h042526b20a689fc88957fa50b,
98'h0f1b8444f704943443a3719ea,
98'h19bea2d03d7c9ff0b188061e4,
98'h022a093294132a7df5ced0b03,
98'h152987dd1304fd11c58f4cec2,
98'h0514109c680535c34a0ba13bb,
98'h0435791eaad6f66deb465197e,
98'h0a0daa3edb54e95d6bc31be32,
98'h1813ee09e7d525b4e958a4e71,
98'h0b39be873370ed95affa44efb,
98'h1805a7424b4730084faaab073,
98'h0f187b91f0f2a8a4a8d335d2a,
98'h1531539e229ce6f97002c90da,
98'h051b722c76f277b3adf38ea5e,
98'h07086522d0fdd988af037a780,
98'h053c62d338f2d7dba6018faae,
98'h000f16045e365527af8bceabb,
98'h0d23bab4074b7f25c7915acb0,
98'h050c9da7d902d6b7451bce767,
98'h011bc0abf7ad658a8783dd17c,
98'h0d1895a2712aeb878e32498d9,
98'h19bd72473ac8bdf3cf90e04a7,
98'h022a8eb9150c825ad5218c0eb,
98'h073410c3280ddf3945cdc444f,
98'h0b00d5e141a8ac618bd07bff1,
98'h0c245e0c88b21d25232a6090b,
98'h0c23693f86f2ce3ca5359ecc7,
98'h0f3489c0a911916fe4c58ddf1,
98'h02381d29301340fd6e1186cc2,
98'h1521ce2c83b6d4c22c92d789a,
98'h0c0cf12359fe6324263628bbb,
98'h0700bd4dc141a7b5c982d511e,
98'h0a2d94e19b3119a222109940e,
98'h05353dd02a558bd36957aba0f,
98'h05091d4b5213c0d96be2b268e,
98'h021f38117e694c9385c737893,
98'h001ce97379f48d99b02221293,
98'h0a28f31d91c078604e845dc34,
98'h0e09b79fd37a5e2426fa5adf7,
98'h151421b36847c991486105710,
98'h0227ea450fe0fb2a0f56fad12,
98'h01129f3e653d7f70a482395bc,
98'h151ffd097fffc8cca99407abc,
98'h19a7dcdc0fbea736b547f1758,
98'h023c29c0384be79cca59a104b,
98'h0e3ffe59bfc2550ccea204573,
98'h0d183d6f7076c59b338094d99,
98'h0419a733f37bcd0baf63c0c2a,
98'h15049d4bc93a1f392de55d0fe,
98'h000f7797decc9c3cc78faf214,
98'h00217bba02d27057e7b704f52,
98'h0a3e39623c5fa198e0bcfb048,
98'h15273d500e58d54771a776bec,
98'h0434bd2029760708a8e004a5e,
98'h0b010dd2421d5bc9eb6ab10a3,
98'h050a670f54df2a6563479a671,
98'h0e0ea5355d52c40f667a645d3,
98'h19a96c1b92c476784ad85a513,
98'h0a123c9ee44cb1b94b1b78a4f,
98'h0f09bee353622bf98b97bb960,
98'h0b3fb3633f414cd8c89afab73,
98'h1989acb253761a9332a0400ef,
98'h0a11e407e3ef52ee8b3ff1d16,
98'h0c012a85c25d49ddeb804dbd9,
98'h0a3b2941b67997ec23979d18f,
98'h0a1cd20b79899262502d304b7,
98'h0f3612f5ac38f731b0e9991b6,
98'h183d8e9f3b2826998edbc289d,
98'h152b4b3916b5b49134d96d4e2,
98'h0a09fa4f53c20bed4af83ff29,
98'h0e11ab50e3694d4a8773018f2,
98'h0f0e6ad7dccf83b5cc5ebe26d,
98'h151d80b17b19b90feaf77ba36,
98'h0b38aea5b167643b940dce705,
98'h18040200480f1b01cf2804b84,
98'h0f2c79d618e361b88804c7408,
98'h0c07f4124fd4e2b0ea03f6e3a,
98'h181d8336fb024755c6f735b0d,
98'h00347eec28e75d1d94c7f2a32,
98'h010c51445881202c4a46f7026,
98'h041b32c3f65eb5bae6635c5c2,
98'h1832b72aa5545043ee9e7a1fb,
98'h071a3cfd745867686f61c1dba,
98'h0b1d01c8fa199d96eedca9197,
98'h151fcd2e7f901d76f14da7d7f,
98'h0c1cd4a9f98c290dd52bfaa95,
98'h180faa1adf4904a8516a3f6de,
98'h0d32b70ba5735781add62bb0c,
98'h0a1ff6b97fd88c2ceca983a35,
98'h0b3b50db36b5aabb327e20b99,
98'h0e32272d245396a5f07c3ee59,
98'h0f1d57b5faa88a738ca16f74c,
98'h0c1d25ccfa4f1b245271788a5,
98'h15252be78a65fd54919b103c4,
98'h0c0da81cdb55362967e2ca4f0,
98'h0a2b256e166151f609d8b7919,
98'h0b11b3d1e35faaa5e8231dd90,
98'h0a1190f6e323b7e18b9c579df,
98'h021453d0e898d2fa6b4d52361,
98'h0d175cddee89c88fcaab49b2d,
98'h0f3e7d2ebcd401f8eee8495b6,
98'h0f2c763018cb006a53049fc9e,
98'h0e222431045e53e169fddda69,
98'h0524d5ab898427c9c4a01e04a,
98'h0f04814d4938ef65a3aa3f5d5,
98'h02173cbcee6dabf6860f5c2cc,
98'h180c8626d93db6a62c213a2cd,
98'h1824a2808956e82aec528f334,
98'h020a8293d51f6834685ee2aae,
98'h0a1550c46aaf5e8f05ca7ab21,
98'h0c3df9993be630108d312bd4d,
98'h0428b1041156e13c72090a6a6,
98'h182ea66b1d79a8ac255fe4902,
98'h0e24c96e099dab3b6d6a13c5d,
98'h021db1707b794be8a5f09d2a6,
98'h0a2269de84cd6984cf65bf564,
98'h0704153bc814541663bbf4d8d,
98'h0d0308e346043402c3c61a549,
98'h0e033393c6420cf6c4c1cf398,
98'h182d50b81a9a768de5115022a,
98'h0d1c9a6cf92b94ba0cb1f1d18,
98'h0c1d5c4afabcc9ee31920bc9b,
98'h0235f8ec2bc80d0251b6898e4,
98'h0c05a437cb52bcddeb7f817b9,
98'h151e4466fc9c3bdfe5d618457,
98'h052d9bcc9b3b8d05b46ea011b,
98'h07390d61323e9cd3a81a4a349,
98'h012afe0695d9cffe6e5dea8d3,
98'h0b2504910a30e1cf25c133814,
98'h0502ca91c5970c50e55579981,
98'h0e22afdb054fe432c2a675b8b,
98'h0e2ef2cc1df8427624dca5037,
98'h0a304f54a08b05d04b09cd509,
98'h0035b6c1ab4c65d74aaed5493,
98'h003ff2423fc401e7cae087263,
98'h072fb2301f6dc5cd9000fd0a7,
98'h021cbc18f9682e2b09a75dff6,
98'h18099984533f66a1aee13a90f,
98'h0d04597dc8842bbacad240098,
98'h153ea6db3d7f4a8d2562214e2,
98'h0129a54593430827d4af7c5a1,
98'h0738b701b176aab8251b2b5b5,
98'h0a057d75caf9ce732e2bd86e7,
98'h0f331674a601203c453fd2fa4,
98'h180ac8435590880ded4d0dac3,
98'h182cfe6199d3bd226b66d4145,
98'h0702a912c549add94c802ee10,
98'h0228c1a5119d1563631315bb0,
98'h0405e579cbd9092664f175c22,
98'h0724a9cc094737e7c3f7bba81,
98'h05387a3cb0eb04b5041af86cf,
98'h022a841415149789ed88dfbc6,
98'h181c6050f8ed6db785cfc6e78,
98'h1802de69c580e411544273821,
98'h0e0081db411aa4cee760f09ec,
98'h0b08f46a51fed33823c6c9aa9,
98'h0700df30c1b83f0b2741f1e8a,
98'h010c4c62589bd9a6e22e478f0,
98'h053ce3d639ea16ee066a09825,
98'h0c1d044efa02d3f64fc9beb10,
98'h1818eb8171eacd689187f6114,
98'h180fcedd5f869fafd280ee3a7,
98'h040ff7165feabadb8de59ba34,
98'h0736a06a2d4da44c48feac7c7,
98'h050a91aad5065017cd21112d9,
98'h073b0c0336274c3406843870a,
98'h051fe582fff4e75e2f58960dc,
98'h183750642e846dc1d14533384,
98'h00160114ec010560d1aeef897,
98'h0c1b14fbf63ba43cab05c19d6,
98'h0b264c040c8b0a3f5095ae4e2,
98'h0f18d6e571b298df25ec5590d,
98'h053b2c273647528b5032dbf12,
98'h040905eed2353bd12ee09fac9,
98'h180bda82d798c845e58f90700,
98'h051fd1957fb3ed2c2be928b23,
98'h012b684b16d8e3dff134efb06,
98'h0c02a604c55195f96601130ac,
98'h010ff3e5dfce1d39c4550eff9,
98'h043a591b349ab13168378447e,
98'h02070de74e01cca5ce3542932,
98'h002f07659e2e44bc840236a34,
98'h043c4e1538967be3e79753088,
98'h0f0aa120d551ca75ef34b27e4,
98'h002718648e2fa72509171ae5b,
98'h0c0f27395e5909246395afe26,
98'h0a2491f9892bee0b0a9a0c177,
98'h0c1d984cfb3add8224d420012,
98'h0432c62a25a2b4a691d61d73c,
98'h021a8da7f51bf337ea755eb42,
98'h19b1fb7b23c63478cdcda037f,
98'h050d88475b086dde4f5e0bfcf,
98'h000138a0c27afd7228057d896,
98'h0407edd8cfc581fec09f0d84c,
98'h0f3af98135e5e6f404f35bf5e,
98'h0010b5b8e153fe127148381d4,
98'h040714304e2170cf08592cf2d,
98'h1981c5f443acc381048a213fd,
98'h0026cdf38dbb9445274ba25d5,
98'h0c340048a8302fa5a378988e3,
98'h00102040604d05064d190bfb9,
98'h1506ff22cdf174c7a8174951a,
98'h051d2dbb7a6ae23388be1cfaa,
98'h1801829fc336e3212fe203fbb,
98'h1804e73949e3d75e86ce19704,
98'h0f378d8c2f3821da287a2fa5f,
98'h1501e0bfc3e9ad880f9bebd99,
98'h0e1332656653580c663ae391f,
98'h053c5682b8b84c212d19a29c7,
98'h0f0d10585a2245c00f7d28a8f,
98'h0b3c61e838fb2a0a2a4bd5861,
98'h04118041e3084cef510de2fc9,
98'h05195e8572a22e9509c6734c4,
98'h013f71af3ec26a824deee3469,
98'h040b7f1e56c702825000770c5,
98'h041df7dcfbf21f51a6b4a0682,
98'h0e3492a82933d102b00405cba,
98'h051586b8eb0c4927cdda18eab,
98'h0424f94889cc78b84c0873f82,
98'h0429dfde9384ebbc437c5c803,
98'h0111c954638b2cb2c5ebb2e6b,
98'h0521af9c8340e9b8c9273d81c,
98'h0a21244f827185732218a6555,
98'h0138d9efb186adb64324aa70b,
98'h0a21bbf0837f01ebacafe1e97,
98'h0b2a778394d6c33de3682f771,
98'h1832871ba52df87c88004eb06,
98'h0b0f82b6df055fc84f581fe60,
98'h0f0fa6e65f67f7f68a85389fc,
98'h19bf3495be5ddbbeeb9de7b73,
98'h0e297b9492d2989bf60744152,
98'h0d0e11dd5c091b79c83f050c2,
98'h181ae99c75c5bd1bca45cb55c,
98'h0e38a7fa315fe843737829ae0,
98'h0403cea247ac43980fe6240f6,
98'h0136fa0a2dc2395342ec048e9,
98'h0d3ca67b394026a24bbe4cd75,
98'h19a59dd98b3c6cd3319f33475,
98'h1988602c50c30e3ac93882ab3,
98'h0f2188e5833370dc2a92db99c,
98'h0d1962eaf2c450d2c4953e707,
98'h0b238d5b8700dc774ff76cef6,
98'h022ec31b1db5644aa4891a74b,
98'h0a1887187117f89d67f909d97,
98'h003ea7533d7dbef4aecc1fed7,
98'h022338a8067cb9372f6f1991f,
98'h0412dd5765af28908227fc77d,
98'h0724d8490985a61dca708179f,
98'h0e2c9f1c192b7b50842a9f99b,
98'h18194ce7f291b41ae9d6069b2,
98'h043487c7293cd4d4b2aac040b,
98'h0e041b21480b0de64b5c5726f,
98'h0a2bb8ae1751372e6583ca41e,
98'h011b0242763fcd29a85f3bf72,
98'h0f032e54c67a99de2dd6b3db0,
98'h150b4947d689a37e455f720cc,
98'h152e45709c846ad54ae53b318,
98'h0a26bbdf0d6d736c8c6cac117,
98'h00356fe6aadf7f7565e50bd2e,
98'h0a3557652a8bd96e4ac53bd70,
98'h0b3e19cbbc15758e6d304c34d,
98'h1818a7e6f16ba4eb91d4e3d68,
98'h0a2cbe6519648462126113349,
98'h051dd5217b97413de8e450b1c,
98'h19b62d282c54bda1702d4597d,
98'h0d0b5f81d6b60eae3182bab26,
98'h0424feb889c7be6cc8f05b8c0,
98'h01278d240f3aab75237b2f495,
98'h020839ecd073d055a4188e265,
98'h19a486d6892f2cbc049f0290a,
98'h073028c9206b7a5d08b4ece4a,
98'h0c0f2515de58479c69e6e8c98,
98'h0d0e5d82dc8281f44a99db2c9,
98'h010d6d0edad86a1e6a6437ddc,
98'h0e3de77e3bd15bfbe6f975cb5,
98'h1529bd9e136bc43b1283d0de8,
98'h0128b85091480dc44a2560764,
98'h1997ac51ef4640dc449c31853,
98'h022f38bf9e717e0f32377b4b8,
98'h183cf47339ec14680ef455da2,
98'h000f9265df0c6ed9c8282db3b,
98'h15270dbf8e38360e27c7004fe,
98'h180dc9c75b9059fde8d7d0f37,
98'h18360d762c2d92610ce788f15,
98'h0c329a13252b54001118e7f5c,
98'h0f3e6437bcc46419cc577b84c,
98'h052fd5971fbdad8ab300b2145,
98'h0200e989c1e001b8893b60c87,
98'h0f212650024d5f3640f83ad09,
98'h0f0aa5205548c82ec45ba1619,
98'h0c1c0aeaf82ca28b8914db53c,
98'h0d3283e1a5070bddd1122b5d9,
98'h003483c3a9017b044c8e63efd,
98'h071c3ce1f85579966a4d7fb1f,
98'h0c236fe806f72f08afdc6d9e1,
98'h0b2566660acbe798c4c6a7bc3,
98'h022b9a159712b0f1e57c537fb,
98'h0e11bae3e3539696e64f92c1e,
98'h050a75b8d4d2f8096c59545eb,
98'h19bb8dffb725e2b106775b709,
98'h0a318beea336498734385c2c2,
98'h153d718ebac664794b59f55d7,
98'h0a3598842b2d71951400f581f,
98'h0e3a0a95b41981efed58c2864,
98'h041056f660b5ec4c3094e3216,
98'h1517164a6e286f85893190d0a,
98'h0701ff7243c3feb550cfe173f,
98'h18309f10a113a11c62b17f89e,
98'h0f0f73d4ded5bfc96e51100b4,
98'h19b9617eb2e4ab038b794ce79,
98'h0f0a1caad4381171332783208,
98'h0f2d61589ae092fe08d08b870,
98'h0d3e7631bcf68985aa837d15a,
98'h182bae93976b913b928d3fedd,
98'h02164d566c9f4ad0ebe5cff3c,
98'h0f3c5a5538bf415dabad6609d,
98'h002bacb59773ce0a31fee6ecb,
98'h00379bf1af24437505e7deaff,
98'h0a39799cb2cf9adbcbd6f7d9a,
98'h0f3325ee26504d036f42451e1,
98'h0e06c1084dbdf0de2d60dcbc6,
98'h0c0aab005579a9f8a6f12c79a,
98'h0419b4a5f367609a8861153e4,
98'h0008930c51212db60de045501,
98'h0e2f57d19eb0548a244a70309,
98'h0f23e02787c3940dcb37eb16f,
98'h0a24dc9989918a15e5b9dd0d5,
98'h043843973093523f64ed99abe,
98'h19afb0ba1f637a960d32e575a,
98'h0a0d62cfdacbd7fc4e44cad40,
98'h15313aa02245b45449364eb30,
98'h0a324c76a49f40666dddbbbd1,
98'h0c23466886bb23892bb463374,
98'h07221d60842f730d04b79a7c7,
98'h010a22e154444b5e42d4641b6,
98'h0d16d592edb3b4f225539b8fe,
98'h07096e86d2f06eecaeb2a2a14,
98'h041f5d427e9ba987667e775ce,
98'h0e289485110eaa3c50aec1b27,
98'h0f3db9d3bb70c3aca7cdcfb05,
98'h0e03f9bb47d7fb4772ab9f601,
98'h180272dcc4e726b30576fd40b,
98'h0217d9b46f9b3af6673a6663f,
98'h040a2721547ef75cac6cc52ab,
98'h0c01d3ae43a406220622479f8,
98'h00325197a4871cd943e976741,
98'h04062795cc459693c92e5b9c3,
98'h070a3e63d44271ca4412ef8a6,
98'h0215a3086b628c0406d32c0b8,
98'h18352fdb2a6065408b5e0bc31,
98'h0f013e52427aa51d30a56546e,
98'h0422b383056a0bbd845ef8dbe,
98'h01386970b0f76876a2632fd02,
98'h0f3227102474a0322c8bf479d,
98'h0e1f09117e20bd9a0ce9b1d09,
98'h05066d674cda74fef30ff1aad,
98'h0a38239030527600647838999,
98'h183ed39d3dab54f50ea2a6642,
98'h07123dfae47bc612b57a8a248,
98'h013a25f7b4755455aae381036,
98'h0012690e64e1ae2a0d6bde935,
98'h0b38f4ebb1f711d2293d05ce1,
98'h052afe3715cd538f4f4c01af7,
98'h07240a1d083c678aa6be14719,
98'h153b0c93363f497b23d81c69f,
98'h0c2c0d6218168c10f2de95839,
98'h198375eec6f0ca17a910a65cc,
98'h0a2759bf8e90a365681d1001a,
98'h180ebbc6dd5bdf7ce62dff494,
98'h15030269c631bff8ad5aa6d0f,
98'h18187c48f0f37cb3a6cd3098a,
98'h0f0c07c6d80d53ad5242fe3f2,
98'h0e319f51232486b509c656dd0,
98'h0d05bc6a4b5310d2ec5589818,
98'h070e336ddc68cd6b0616334f5,
98'h0b325a1a24bf3b2b28ddc0363,
98'h1999fadaf3e4f4ae0bfc65515,
98'h0c22c6cb05bc68e6b35fbbe23,
98'h0120a885017a4d46a477cbec7,
98'h021289a2e537b3a6a0a6bd72f,
98'h0e06cd0a4da59dee09d28f526,
98'h1804eff549d8597c66eb1abe1,
98'h000073b740f3dc4e2877525c7,
98'h18086247d0fbcde8203d14016,
98'h0d226f8904c5d5feca410c0c0,
98'h0d34e94fa9c73adbc47a1161f,
98'h041b582c768bc9894dbf090ad,
98'h0a2ae2f195cf71b74ea9c86d6,
98'h041136fee251ef66e7fe952a3,
98'h0a06e7434dc84c4cc998c9997,
98'h0c10e40c61e6f2ff85f3cce40,
98'h19afdd889f9c7ddc6b7df5c2f,
98'h052c131298155bae6e5316d94,
98'h0a14413768bed417a7505bb04,
98'h0013107ee618e5ba6cb4c553c,
98'h001b96f47735e81f298afd8e5,
98'h04272e6d8e68cb5d8dd45fc4e,
98'h0001119442133f8464a3fe72c,
98'h0032e1ac25dffdc0e08514463,
98'h0b3c671c38f6dd47a984b7db4,
98'h19a48eb7093c4dfcb10cd118f,
98'h0b0dd5c1dbb042da28b8372cf,
98'h0f1906bc721d861ae9af86270,
98'h023258e924bde11db04da335d,
98'h1832b497a55d7213e9bc0e81b,
98'h00350e282a1bf962ef6409aae,
98'h182a79d694c9d8d04a9441e2c,
98'h0002ca434583ee69cb3d14a9b,
98'h0a373bb6ae79652a2161ae2b4,
98'h0414de2f69ad05640e2c28383,
98'h0b19202472647ee98b7078e4d,
98'h0a380c11b00f96f34f5f67c37,
98'h0d057abccadb13c8ee91e8c13,
98'h0b24ac3f095bb027e5f823a17,
98'h0d2069cc80e0506f05201719c,
98'h0f0d023cda042382c3802e8ee,
98'h0a212351026549768a44496fe,
98'h0d36c1bfadaf09f503219b31e,
98'h182df1f79bcb94684eb972ed2,
98'h1824c3ac898cb3e04cfe6197f,
98'h042ce21c99c8d0bcc86c5de33,
98'h0105eb194bc60a14477d6cb65,
98'h04361ecdac3420dca332fd4b6,
98'h0e0e3a495c635ed28c1a8fea9,
98'h0d04fec6c9f693222a9c6646f,
98'h198f17b35e3caecd25bee47a4,
98'h0c34c17629877ad54df2f1a02,
98'h1513c2fae7b45223ad6f0f12d,
98'h0a05fbf7cbcdb92fcf320547a,
98'h0236f9f5aded1d678574ed49e,
98'h0b19b619736ef6598c0905d74,
98'h0216cda96d9cf29a6fa22b1cb,
98'h0a3f3757be45ca6ccbecf010f,
98'h053ba749b74cc22c522140711,
98'h0e2183df0327d6718f221a5d7,
98'h18377d3c2ec6fbfe445256942,
98'h1511898de314cd61f1bf9e4e9,
98'h15323815a46570620e0995bbf,
98'h0e19fcf073d76d256e65ea1de,
98'h0108479bd09fa118707c5a857,
98'h0139e64333d167966469fa2d1,
98'h0c1067c360ea82518d42d3766,
98'h0f12de73e59b3b7ceb3eba853,
98'h020d95b05b2aabaf8d2b867c3,
98'h0f07fc1f4fd0fd92e74e1057f,
98'h040234b8c469f94307b63e6c9,
98'h0c3a709234d51180621b0b7ef,
98'h0a096361d2f19c8d3043e084a,
98'h0100d4c9c181d2dec73ebffbc,
98'h0b0b805f57199d7ee0a0a9ea2,
98'h002626730c732e37288947779,
98'h1512df97e58ecb78c326552a9,
98'h0f2d74eb1ac12a02cea86ac42,
98'h0d35af1eab401e4bca7ba7bb7,
98'h15073e3ece745fa9ae1d735a9,
98'h013a0c3a34148739e8dee77a2,
98'h05157c2b6aed64860d53a4dd0,
98'h0d09485ed2ba31f2ac00b82c5,
98'h0f0b611d56e822e007f0de946,
98'h0f375e31ae903598697ce0ff5,
98'h0125c5320bb422f1af71e4f28,
98'h15139687e71bb5bb63367a08f,
98'h0d29433692aac3e28f0bd310d,
98'h02275d660ea9735c87f501c64,
98'h000305a7c61c64cce4343430a,
98'h0238470130accded8187da9d3,
98'h199943b2f29d7db8ecb9453ba,
98'h199244bee49d344ef30db05af,
98'h0c086e3450cca89fcf8bde437,
98'h040f0a33de0305d1c73545b50,
98'h0f3a0cb9b41a9a6ae88484016,
98'h153fa224bf54e336f0d529c92,
98'h0f324a7f248d0bf255252156e,
98'h010d3386da766faf2cefd59c5,
98'h182133730265930006e0e8cd8,
98'h0415f67f6bd981dce6a1b19cc,
98'h0434a13129456b4ccbfbde171,
98'h023b5962b6b2c4cf2b5e831f7,
98'h0c17d8076f972f816e3b878c7,
98'h070655b64ca2c9078eebc1e23,
98'h183dd3f23bb78236a4ea47af7,
98'h0436f52f2de4857814fd558a3,
98'h0203459e4685a6f64c86dea9c,
98'h0e0406b24802488142223b252,
98'h0c253f690a750b38a58193cce,
98'h0d000354c00218f345a692a87,
98'h183992603328bf67034087120,
98'h1808235b506a871012d89471c,
98'h0105db3fcb91dfda6a1caa9ad,
98'h0b12a33ae570ed882325eec69,
98'h18023f74c479eddbac20e430c,
98'h072138988252227ce71f0b542,
98'h0204da1cc99218a3e25cd6c56,
98'h0f0cb749d946987ec2e5bcb03,
98'h0502d9044590765bea14d3f22,
98'h070ee652ddf2ef8f22a4d3d81,
98'h180449a848942d1ce94075788,
98'h0a1f84e97f25f61f08261db15,
98'h011796366f398befb2515ec21,
98'h0e297f7192e51a0f0c1448898,
98'h1981b28ac37713cda843a6602,
98'h180d5481dab849b1273e31962,
98'h0417f932efcc709fccb1678cc,
98'h0d15a9ddeb5644c56cf91a74a,
98'h0b20b86b817c623e2e1afba8d,
98'h0433117aa6025d7d432746aa7,
98'h19876f224efa95732a8d5bbdf,
98'h0c03fe7dc7dca9796a2081256,
98'h0121b9f383666cf684f829fdd,
98'h0a1dea3cfbd5a2cae12209ba8,
98'h0531f02ca3dbba72717ce341f,
98'h0b3ca93b396638f28a436aa7c,
98'h0d0470ca48d2677ef128b88b6,
98'h0a2cf02f19dd51e1e575b6125,
98'h0d349f79a9360ea5290290844,
98'h053708fd2e03baf9cd9aab87b,
98'h07169197ed0e845eccceb0fdb,
98'h013eb7ba3d478a0acd09457da,
98'h18326b3124c250144fa190713,
98'h003d4fabba8fee56cf3d2ed15,
98'h072e6c039cec151e0eb34f809,
98'h0e2af84695ca718dc906a0486,
98'h0234ac7c296bebc688fd5a751,
98'h001c222f7872a8d12ae82610a,
98'h01118ab6e30daa45ce23b2c02,
98'h0f082c3b504555b24907cd3f2,
98'h0237c7812f8d1dc4c7d3607b6,
98'h0d1e386ffc7ff731ac7139517,
98'h198753584eb1335cb2678be86,
98'h0c3d31013a7dcac0aa0e21ad4,
98'h0c23cb6907a7111691aebef07,
98'h0c13fd54e7f33d4024f2b71fe,
98'h0217a690ef761eebad01cea54,
98'h0b1ee6ff7df8cc00ac63715f2,
98'h0f31125c2215ffc4f245ecc00,
98'h18272ec60e4655c3cc51c4884,
98'h153580082b1f7a7a699b61227,
98'h1819d19e73afdbba90153ea0a,
98'h0738e181b1c152d652f26b563,
98'h19ba7dacb4e4b2858e3e8d15f,
98'h02159665eb121290f3a7cc0c8,
98'h1527b7460f6223360b49ea3db,
98'h01320901a407c2534922769f0,
98'h02152df06a7a7c4d294e72d53,
98'h0c30fb52a1ce92b6cb23ea8f6,
98'h0411415ee28192bb4b7fe3825,
98'h0b1984057327754409a4b5068,
98'h041ab678755fb2e26f903e525,
98'h0233bb762767a5748e5e9a56b,
98'h0f3b9c50373c0192aa66d83aa,
98'h0c0718b2ce2221b1119de778b,
98'h0b0e612cdcdf4d0d668a4e98f,
98'h18177e786ef4145229fb6b8e9,
98'h1982178244204e0311c2e4b2a,
98'h0e2df8331bdd2ca1e76899615,
98'h0422eaf605da5895ea82c9354,
98'h002a2701147ce7d7a27f50e30,
98'h0b1bc55d779f7d55e529c3b63,
98'h0b095eaed2bdca1db0aed0acd,
98'h181623bc6c471a444771ca332,
98'h010072b8c0e7878c91174f802,
98'h010d1b48da29dbd20079fe915,
98'h0035334caa411d2dc6cdbdc6b,
98'h02188e67710c2de0ca9d941e9,
98'h00149a47691bd9f9ecc92f120,
98'h0e2591ad0b281cc00a4c1d105,
98'h0b32a835255057d9e6536b9b4,
98'h180100df4237a632ac20c003c,
98'h0010f15461e664a6068e29c48,
98'h180943f252907a68687dd57e9,
98'h1998da90f190db296aa66f96b,
98'h040c440bd8922d0272ca6d6e9,
98'h000686884d166c1ae7279c439,
98'h0a0690804d17d611e3473ca8d,
98'h0731728722f0572425c799a49,
98'h1528b3d4914e2317ca88726ad,
98'h040fc38adf9813dee99db5bb1,
98'h0f37b8beaf7ed80528e9f5da7,
98'h0a01434042acead30fada430f,
98'h0e0ddf22db92c03ae32b8b84d,
98'h001f0d047e0a7e7aca6827d77,
98'h0c308116213b0f8a2f8a62dfc,
98'h053ceae439d9443e6b5ae4281,
98'h072027dd806333338fc58bc8a,
98'h0539629cb2d1ed76e1e0d6c44,
98'h0537d0ee2fbc12e8ae02d404e,
98'h0f29729a92dcc06ced3cf8f5b,
98'h022062ed00e1c1ca88818cc1e,
98'h001cfefb79e5e15980c0892de,
98'h020d52af5a8c9f69ce80b8153,
98'h1828ee8b91ef8b6687267c864,
98'h152778390eeee8c68a861e7c8,
98'h1993f7c967db39ad6905983fe,
98'h0a3b13c0b60fb953d05bcc5db,
98'h0d331ddfa612c034f012b3451,
98'h0c2e02aa1c247bf10cd177852,
98'h0c32ddada5aa54f78a149fa6c,
98'h1833248b2659cbefec774ca94,
98'h073a0abeb40488decfa33c1ec,
98'h021ff027ffecc6110ecfa4e75,
98'h01035c50c6b130c2b0832d8e3,
98'h0d3938763265c98581ed2344e,
98'h043aaa5035703e6c2fe7c07ee,
98'h003c219a3875a8eeae6aba2f1,
98'h011ada5af5b18994ae2c72a23,
98'h199845e9f0a64b5d0db318fbe,
98'h0c397cbcb2da88e5f28fa451b,
98'h0a000ae9c03fbd522fc50168a,
98'h051d19737a0afaf7428ff20f0,
98'h1524264e8872b1beafca051aa,
98'h182b2d2b96497f52c765b6035,
98'h0e1f52fdfe8973034b9d2b1f9,
98'h19aad64295b11f70b32a31804,
98'h0407360bce5043f1ebd6fd6cd,
98'h0d0931c55268c7bb0495de7f7,
98'h000773be4ed630ca67dc7e601,
98'h0f3c6870b8ddb08ae3b769223,
98'h041bf48a77d7503ef206863ee,
98'h18126bb1e4e9b7278efcd1325,
98'h0e2f5a139e91746f6f3f08b65,
98'h072862a590fea6cbab3033a0c,
98'h0512a430e5744bed2609c25c5,
98'h1837c7192f9f71a06aa1bc078,
98'h0f3305e6260df2b9d1f5ce2e6,
98'h0c1632896c6059bd0d503e27f,
98'h1522ea6805c4f3454e1da3119,
98'h1834db2329970a2c66b9f76b5,
98'h0e3b2a1d3660b7719072f953e,
98'h0b1cc0c3f9939fe5f126f863a,
98'h02096f98d2d1698f712c182a7,
98'h0b1489f8692ba2d38536b64a1,
98'h0530cca0a198455fed100b32f,
98'h0b0d10fd5a0feecec9b244802,
98'h0b117f29e2e1591309473ff30,
98'h0521a0bf83568c9f6b7cb60f3,
98'h0d3ce65939cfb64b421e0b57c,
98'h1828e1dc91d17afef1c327291,
98'h0b2aa783956d13188a7e9736e,
98'h070377a1c6fb6796a825eea70,
98'h0d14032e681ddafce37fb7ce2,
98'h0d054d0bcab357ff2d4c778ad,
98'h070a5a0e54aaafe805ee2942c,
98'h0b0691c6cd3042c1a6ed427d9,
98'h0a0de2085be05b3b860db5222,
98'h0a19673172c59857497b8f50f,
98'h0a198b31f3372ec92f37bfe22,
98'h19913d56e241bc284f542e7ec,
98'h0d0914cf5222d5d08ef4be5fc,
98'h0c38dff5319f6d8ee7cafaa7f,
98'h052e52559c9b96046f7613610,
98'h01043379487320d2a8727a168,
98'h0f1aa06af5620083825dd5130,
98'h0d3aa200356d482e111f283b9,
98'h071189e2e32e12e090a9fa8b8,
98'h19873856ce7a8cc92a8fe730d,
98'h0d099cc2d32ac81c0a0071480,
98'h000b72f9d6faf7bd280d1937b,
98'h0a106f4060cf19a6c5c19aadc,
98'h0e01bb16c3790b132ab7e239c,
98'h1816d4bfed957062645eb18a8,
98'h042c938a1939cac4316b11489,
98'h011a42d6f482859f475997939,
98'h0c3f75e13eeeb5b88d67321d8,
98'h01106649e0dcb41e72cb8ae66,
98'h011e5f597c82aecac87b469a1,
98'h0229e80d93e4b9108f6843890,
98'h0e010ddec22ad5c20583a8478,
98'h0531624822d0e517e40af8e83,
98'h0136ed0f2dd450596a0091d80,
98'h003b854db73bbd442bc2cf5a2,
98'h0d38b33731780337adddd0a47,
98'h000d6ca35ae70c170fac2d9bb,
98'h19a4ae53894d3af746bd1e2e9,
98'h050e23fe5c64628188bc7a52b,
98'h0432c11225844520c85ca19ff,
98'h00085c4350a408e48a6dc18cb,
98'h021d0fcf7a21f92d042b1949f,
98'h15315087a29b6010ef0fc23f1,
98'h072a5d98148531854df32c262,
98'h0119db0ff3a3b24706ebe3c75,
98'h043719292e0f3482cd2f6355b,
98'h0d1eba51fd6274398c91936af,
98'h070a19f0d4180d6df2a04ba2d,
98'h0e1d05f17a3bf60826c889d7b,
98'h01320d0a2407d58052163efe6,
98'h181fd3c47f818444494e78a29,
98'h15189243f11dece275e856022,
98'h0a2c0ccf983bf8eeb18d9fc99,
98'h0228091a101f23ad689a016f9,
98'h053f72483ee3bc788491cb31e,
98'h02110db9e213d2ea7108cbb02,
98'h1807d292cf8736c2c90938291,
98'h152ca600196ee59209e3c2556,
98'h05076e444ed0b01eeba6e2e48,
98'h0d281e7a9026d18d84f60798d,
98'h0c0b8d22570ca24cc753bc020,
98'h0c179765ef3980b6a8c60bdbc,
98'h0f0a4321d481797e4ed446072,
98'h0c3c41ae388429d548e2ef280,
98'h042c656698d9c55471301ae0d,
98'h043b4bf1b68819a347418aaec,
98'h0538af473151d9dfeeb0d9653,
98'h19b27f7ca4e56bc88da2a249c,
98'h020517484a09e0a1cfa5fad14,
98'h0a078d4c4f04b3df4303bdfa8,
98'h0503541dc68d598b4643104ae,
98'h183f0b0dbe18966fe2e42b6a4,
98'h0d2d91ae1b110bfd7595e85f6,
98'h1998201df05051f36a0fa76ae,
98'h0c08560d509867c8727a1c845,
98'h0d19e28973c437d247282f757,
98'h0b1e9680fd23562e10378696e,
98'h022f640d9ed51566f2107b2bb,
98'h000cfc7d59f57adf28411e5d2,
98'h051f6f17fee78cf886809dd72,
98'h19a15aa802b7e4fcb101bf041,
98'h0f1cf3c4f9d45ec267164fe93,
98'h0d0351d646a63017923c54a1d,
98'h0d1d24e17a56a1eb64ea607b7,
98'h0f0b260cd668153111dcf1b33,
98'h041044ea60b0ed8d295ccecf7,
98'h181bc37ff7a86bba09304c9de,
98'h0f0a230d547271b133f10bce7,
98'h0b04f39549ea9a9308df252fa,
98'h00174826eeb50050253be38a1,
98'h0d22c1e2058f790e4bb3121dc,
98'h002bd3c4179d065364ac8ebc1,
98'h041f112b7e2a9feb05f23685e,
98'h04090921d2147492f0926c459,
98'h002a606514f92a5ba5875f6d3,
98'h19a68c2d8d2998d88548e2b03,
98'h0d30bfb5a17ae70129b409418,
98'h041c4e83f8aae6dd0baae9adb,
98'h053ff5713fdef8ebef31cd583,
98'h013a2c71b448b149d147bb974,
98'h0d03d31cc7a4e89c0d60b76ed,
98'h182a39f49475d2b7252a2eee3,
98'h0d2dba6d9b432504cb28032af,
98'h0f2abfb8957046aeaa1c37dc9,
98'h0f0c5248d893f485e926c199d,
98'h071ce81bf9cab2a949e811b3b,
98'h18086bc350f9d5efb039e6b14,
98'h02151c2aea3fdf0faa40906cc,
98'h182c1721981c5184eb153ecea,
98'h010a10a25409203acc121a29a,
98'h0b08e8d951ce39f4c544cc374,
98'h0a2f82ef1f20af740735c8b38,
98'h02026e8f44de5d616a540c98c,
98'h0539a62f3348f3f441b832fc3,
98'h0231d4182383a65b4e20a688d,
98'h0436402eaca1bbe4096d5e9cd,
98'h1507b8794f45ace3cc35ff04a,
98'h0118766af0c4655d491359574,
98'h0a0132e7c272b76bac7736f20,
98'h0b044b10c88ff768431cfa94e,
98'h013507c82a242bd384e5109e4,
98'h0216c9fd6dbe2afe2ad64ce6e,
98'h0b2e0db01c02706dcbf53d3ee,
98'h0b17e5bd6fca640849cc1f877,
98'h0737c2642fa93cf98eb892716,
98'h0e33048e26239a5e8db83fd76,
98'h05320fd9243d5ba9ad15a7bb2,
98'h0d033d5cc65232cbea5bdae0b,
98'h0531413422b4da1da4d55c0a3,
98'h0f3044c620aac80709f986d47,
98'h0e1f27cb7e42aa674bf6c3334,
98'h0e090a175216e3baf318748ca,
98'h0f027021c4c6b4074807fb749,
98'h1839044cb22ca77f04f2490a4,
98'h0e0126edc25354ee72996af2e,
98'h00252f140a7e65dda4151ef71,
98'h04236e1386c9527e42a8e53c7,
98'h0e2db7ca1b7b2b4f22bb30247,
98'h0c0b61a8d6fb3a872a6a38c65,
98'h0a015a7bc2a9373c88c1a70c0,
98'h0d072cf24e79344b232aa46e1,
98'h0d1f6ee67ef364fea6e0184f6,
98'h0d124f656496417a7304b4f94,
98'h0c15a576eb7284df2c6a2437f,
98'h010b11a5d627ef358de20a958,
98'h003674492ccba51645ccc036d,
98'h04112a89e271770eab408657d,
98'h0d35342baa6c4acd09a0a8662,
98'h0e329416251b50066de85fbe2,
98'h0004ed9ac9dd9b1d6cd379072,
98'h023b907fb7082f8d4278a22e1,
98'h0d06d5c3cd97740f6e50f0033,
98'h19aedf2b1d887a84c6a79274d,
98'h0d057b834aec759c0dcdd66bf,
98'h0c1b21adf65d263d65fc7c47d,
98'h19a9a4669357faad709e11fad,
98'h183270cca4eb09780b4067c50,
98'h0b05d9aacba7021a8f475e912,
98'h0b39217cb26f9d6705ab36f15,
98'h0a05a53c4b6507ae8f6a2fb8e,
98'h1510b9e361782eaa255aab3ab,
98'h003d7eb83ae5cd210da23a236,
98'h07141654e80c7e52cec8d2f64,
98'h0d08686c50f5131babc82529e,
98'h0229be56936dd2e1877f5ee20,
98'h18103c55606542370565e44e0,
98'h1521699d02fb7947ae1d5fa31,
98'h150da91fdb6603fc860738b93,
98'h0b21b50e837db5e6ac1ceb471,
98'h0a3cdf28b9bbcbe523a7dabd5,
98'h0e1b07bef608258f50fe2ac37,
98'h0f33ed7d27e150599108cb538,
98'h0f24a7f309548e81edc54f75a,
98'h0737cedaaf8bf3b2c61e4d9d4,
98'h01190020f227216f8db0f0a35,
98'h199d26adfa7c1d3a2cd008641,
98'h19b613ecac3d2a7a350650fa0,
98'h0f31ae13a3728228317ccf99b,
98'h0f37252bae7732322ca90c0ef,
98'h199b50d976935ea66f6b95d77,
98'h0f0c88e2d91f8e98f40babdff,
98'h0109fa7b53f09ecd2a0b05def,
98'h0506ac474d5e641ee53ea6522,
98'h0a0913275223f7a6049944199,
98'h073949bdb29c16a5670b42b35,
98'h042dacb99b51f02a6e755818c,
98'h000bcddbd7832a7cc7dfe7390,
98'h010e5fbfdc9eda4265e3be162,
98'h071bec65f7c29567476b4e809,
98'h0b21d876838ebbc6cfb7a0734,
98'h05076550cee17f9483ac250f5,
98'h051113cb62392781a4fa39395,
98'h1821f9c203e574a689d28ed34,
98'h053a4c5ab4aa062b0701db9a2,
98'h150c910ed93c04ae2e7914a16,
98'h18119771e3384f6cab92256f4,
98'h02128dbb6508d52c4ed279b7a,
98'h0c3c320d384bb2df49c6d8b9e,
98'h0222527d04a922119121f93b1,
98'h01337ddaa6fa310ba1b2dd23a,
98'h0f25f7390bedaebf0a0b6bb99,
98'h0d2cae369956a46b66c4e97e0,
98'h18312e04a27c2706a9a0d4a88,
98'h0c32252ea4793a66aeab5542d,
98'h1529582412b8f0282c2ad7e55,
98'h010b807f573adc5729f892131,
98'h003ccb0cb98a69d546119735a,
98'h19815695428c88854e71cd387,
98'h002e45639cb69f2f270377c6a,
98'h0c39a38db3439b2a47393924b,
98'h002993fd930c67c64fdf4fadf,
98'h1519e63673e4076f04cd7ef0f,
98'h0c0666dfccf8f89b323f7b695,
98'h0c0bed0bd7e1806d863fd7dec,
98'h050e563f5c9ae52068fb5b5e5,
98'h0432533a2480922d486a4ed7f,
98'h198b1780d6139035ea2cb959d,
98'h0b09ada05370aaa82be7a9edb,
98'h0711e239e3c80d2c479e96122,
98'h0c2367c906e812c70ab67bd98,
98'h1831052e223270c5a4c2dea40,
98'h001750f36ebad7632e98dd7cf,
98'h0214ab54e95492326bb48a15a,
98'h0c38d90ab195a244eada4f61d,
98'h1527d0d08f8d3c134f739ed3e,
98'h150cfdad59f58325292d4338f,
98'h0c2667f80cc0cd79cbc0a034a,
98'h152de7271be5a8ae0639cd5c7,
98'h0c05ae504b764ae6ac44e3f54,
98'h15393575b27c0977a5defe4dc,
98'h0f07b18d4f79df4b31ed4fbb5,
98'h0115fd466bfdfd0b27a064362,
98'h0c3f04943e05cd07cb44fe946,
98'h0f0f74f55ec5c4e152913466f,
98'h0b37a47a2f62ceee0b754e75a,
98'h0d31518fa2b20563aea69cda0,
98'h002a0d849420e93e8bf8d5bcd,
98'h0a02d3d345982eeb6512bdb0c,
98'h180d8028db39aaab23e6c0afb,
98'h0e2d852c1b22d6c00cd1cab50,
98'h0c0e760a5cdcdd53ea5416fb0,
98'h0c0ca4b85975001c2a3ad4d79,
98'h181e46ff7c98a7c9e96069352,
98'h01124443e49b5528f52dbbb25,
98'h0500fe0cc1fe1e0e296b665b3,
98'h181f154bfe044ffdc1bfc706c,
98'h042e5e669c934291f588d9526,
98'h1999e5fdf3e853a48830683e2,
98'h010b1873d613773673608e689,
98'h0b03ce3647bab51625c7a3ea9,
98'h0e2f2ec71e6f5e4b84afa0d32,
98'h0a360c82ac2cb43c0b27a344a,
98'h001e8b277d2d2b940d98b02fa,
98'h0e26931f8d3b64ef2f52edaed,
98'h0408c38851ba653fa6d87e03b,
98'h000044fa40b187f7a570ca320,
98'h15150f0fea3014efa02c733c8,
98'h020be2af57f6540f2fd148ffe,
98'h022f6b121efa68b526808dafa,
98'h0d16a78c6d722edf284a74f1d,
98'h153bf014b7c4c4114ea2359ae,
98'h0c33968e270255ffd3402d097,
98'h198556cccabb40f4accd7b237,
98'h0b24776108e477fa091025f06,
98'h022bad1e9762a0c005023bd6c,
98'h19a783638f333d47a6639377a,
98'h07083b205077ad45aa36b02ad,
98'h1996c2a16dbcc150a5dffa198,
98'h0c2b9815973709c531d4e0fc8,
98'h053618d7ac2bfb6f08d8a876b,
98'h0b0aef7455de73f0ec588511a,
98'h073d0273ba2e17eb083a58d95,
98'h182175e102e874e8105ac697a,
98'h07190192f22cc0fe86c27ab24,
98'h0d3b0e313633823d2e5170a45,
98'h0215bb016b6657d190dba41b9,
98'h0c0d1e695a358ef0ab5f04b4b,
98'h0d07c33c4f9d1d7de990ab568,
98'h153294bea50d0c734729382e9,
98'h07071b714e064c0bce8fe84c7,
98'h15101c9660305ba6a54359df4,
98'h18365e7cac921f74ed501e0f4,
98'h181583856b2caddb91321f7c6,
98'h0c039debc715cea170d08c583,
98'h15014e50429555d2e4c65b235,
98'h19bfeefbbfd0746b65e5a908d,
98'h053b7dec36f488bd366418d9c,
98'h011aa7997573e89aaf0c01aa5,
98'h050c847ed93e8f3c2da3a40d0,
98'h0c3d4b61ba8a88e9c792c4eec,
98'h0c256a5c0af86660b1b1f512d,
98'h183528a1aa42f20045c7742f3,
98'h0a1e2309fc72d0abb09e06a87,
98'h0707a5564f5aa877f1a43ced6,
98'h0b3f123cbe2ad70e059893739,
98'h043e3c2cbc50b1d9725a7a52a,
98'h0a1ac0d9f590b9e97023bb818,
98'h0f2729818e791d9dafeadeb0d,
98'h0a2cc1f619a6520d076811c7d,
98'h1537c862afba7e2da8f4c500c,
98'h0022c7d60595e1bbf13c91a41,
98'h0e2d9f8b9b2e51e3016e2a648,
98'h0724e8f009d255a66a56fc5ba,
98'h0f3b1e6b360d5c06443dcfa5a,
98'h022214e78401f5ecd1521e9c5,
98'h153d0a1cba00edd0c18902b51,
98'h0a15b992eb64872093cf7dfb5,
98'h15259a6e0b221f6a8d5e902cd,
98'h0d2b97f61715db436811ee762,
98'h043a46dcb49ff8ede9105cce6,
98'h0d16c946edbdd2c52e368ff2a,
98'h0531439422b58b62aeb527030,
98'h0c20f3e901eecd8709f9b3bdb,
98'h0d2bae729748f9c2c383f05c0,
98'h1526b0728d638bdb091d2a0d5,
98'h15396c0532fc71f628a28f136,
98'h07261ea88c3d7f81320d777ed,
98'h0e03b488476a15d704d8e78a7,
98'h1834aa8029548caae55b7297d,
98'h0f2b50e896b3d42db0624dcac,
98'h0e21011d02193af8e977c9459,
98'h051787c46f0031b3c40e8f058,
98'h0f3635d5ac7a567c2d05ee5e0,
98'h0a22ba67056d02110eec23147,
98'h1985172eca2f00b603e3ef1e0,
98'h1501b1cec37110dfa8ed05f93,
98'h0f08b3dc51763197a61cb0aba,
98'h02329ba82515baa8681fb95d0,
98'h182b0fc4960ca881c9d215942,
98'h0f30b750216175e38b8dee119,
98'h0a1f08fbfe0a4d44cc248b4ce,
98'h0f19b2d3f37c4bfab20a55902,
98'h18346cc728c80122d0a57fb3a,
98'h0b21b7f003474247503f1b7a7,
98'h073b3c9bb65edfcbe39a3e8dd,
98'h05232912064fb3114f668719e,
98'h053b231eb641f06142dcb708d,
98'h05070e574e379692aedf44dff,
98'h19b41924a823467404cfa93a8,
98'h0233328ba65bbbf3f075d7e62,
98'h070d3ab35a459305ca23bb9fe,
98'h011af02cf5f0f24da854b36e4,
98'h0406cbfe4d8b2586cdc2f89ea,
98'h0f3fae67bf4121a9c4647c614,
98'h19b46e6ba8c35cd7d3a034045,
98'h0a1e0e197c215400909df2d0d,
98'h04348590a927884a918fd8867,
98'h0e34c6cea9a9ae3b8b570376c,
98'h0009cc31d3a8389f8df79d428,
98'h150233c44468593304ec81345,
98'h022c1943981c0108665aa33dd,
98'h0e0590e84b385ab1269206930,
98'h0a1554ec6a90a825e64f7ae66,
98'h0700e7d641d55e6ded297f449,
98'h0e3f9d7fbf2fc908023591911,
98'h0428acdc11756f12335bd9a1e,
98'h0b399c833317e430e56786fb9,
98'h001e0bf77c219f378f94602d0,
98'h0f260bac0c3ae0912f0feacbb,
98'h1980e5d341f6a26726d83b0f5,
98'h182b69df16c2fc8a46dde20ea,
98'h19967cce6ce656198bbb999a5,
98'h1988e031d1ef2eec119f34b9f,
98'h0f31d1f523833ab84ade03c77,
98'h0d3556e82a87f7f94cad432b5,
98'h183ab204b54edc9b4def53b85,
98'h071dba77fb7da261336263a7f,
98'h1820726980f42d0cb0a6d7364,
98'h01077085cef0f445a64527dd9,
98'h02355e41aa86cb44c3fe1932e,
98'h0d0bfce6d7d75037eb2f0a619,
98'h001fd3597f903d6ce938d347b,
98'h0a12d69fe59b46386fec04319,
98'h0f3e0f2d3c24199d8beb87361,
98'h0f1e6ce67cca94b852d88a32a,
98'h0109abeb53641ee092fa4067a,
98'h01315c1ea2929998651b72b2f,
98'h0f37cd6faf8d3e2ec8f0fd6dc,
98'h0f00d2dec1bc332a2fb142e79,
98'h0402fe47c5d69370e42f41824,
98'h199926eaf248112e4276646e3,
98'h183bbcb0b75b4e7f72f84e064,
98'h0f099a37d33c75d633e5c2cc0,
98'h0d2cb79719788c24289184038,
98'h0a1c4feaf8a566c209a950eed,
98'h150fbb98df781f17b0b06dab3,
98'h050f7159def84e03ad21f6ac2,
98'h02005001c09149036901efd76,
98'h19b48308293c0b1ba0a466415,
98'h010903cf5238637fb0bc2388f,
98'h198ae9ac55c673fac4d059d3c,
98'h05186aaef0e679160bd45769c,
98'h041a9f2a75104602ed7fb8f13,
98'h051ac9fcf5b1ce3fae4ab94b5,
98'h0704179748108703eeb3260f2,
98'h19a575c60ac05a6543c527a6d,
98'h072a56389480563fc919740ad,
98'h0210ddc8e18d30df46eaab1e1,
98'h050c3283d8582d66e8e783aa0,
98'h0b0e4a715ca9d9f7875917fab,
98'h0011cd1c6387919a49ee091a3,
98'h153649dbac949be6e8e657ada,
98'h0c0334d84658346b7072b970a,
98'h153cccd639acb3d58496da50f,
98'h180d3bbcda5d84daf3ba602ae,
98'h0427f3dd0ffd7eddac9ab025f,
98'h0a297bfe12c1b059c5095caeb,
98'h19968c1e6d099307c73acb15f,
98'h0d2e8d019d3113c931a807c98,
98'h0e133c75e66ec84c8a97e832b,
98'h19bd685c3ad51c79ed2081309,
98'h0421627102ec31959524a1358,
98'h0f30fed321ff992ca1c36501a,
98'h04209f4d010305bb4c4c25fff,
98'h0124fd5b09d77b13e148e9421,
98'h011414f6e81b788762bf1e1bc,
98'h0718c219f18806ceca4be35f9,
98'h0f0a530ad48683b1ce28323a2,
98'h012381630723756f08e435af2,
98'h0a12f3d6e5e59fe40211bdb48,
98'h0b1e9abd7d1a05766bfe24eeb,
98'h051ee957fdf16db7b20e280cf,
98'h0d1b1ddbf6167bd470c415c3e,
98'h01187a3a70c84eb550cc666c1,
98'h0d277fa50ec114eb4c78323be,
98'h002feedb1fddee55e6fa25241,
98'h021a7f2d74d9e58be803774c4,
98'h0b09ee47d3d4bb026dbd192e5,
98'h0c083ab9d04babf647b7aa529,
98'h0d2c8b3d193a4f132714f9ac0,
98'h003674bf2cc810dc4999b6941,
98'h19b80128300fc9d2cb3fa166d,
98'h199508e36a2e585e9271f2beb,
98'h0528212610771878b0f0d8507,
98'h0b2f90fa1f2d830e8567ce67b,
98'h070b6f03d6ce2f2eca9745022,
98'h0a3d3a093a42deed4776678ca,
98'h0e0cee3dd9f1320db120063d9,
98'h0723c94587a6086b09ff8812e,
98'h001d9f01fb0c8e1ec3b2746c2,
98'h0432d11425a35b698eca8b482,
98'h003aab2c3558025aea758b1f6,
98'h198c160a5815d4396d64ab61c,
98'h0a3d434a3a8398aacc687a90f,
98'h199e23ec7c61609b913036fd3,
98'h00112b99624f8ee7557fe121f,
98'h020612af4c3ea0c128982ea02,
98'h071ef905fdf82fda23912cdc2,
98'h041d7b78fad9184b7145ca380,
98'h0526fe2d0dce9c3bcfbda4f11,
98'h19a99d9d1330cf4aa4bd669a3,
98'h19b9e85c33c783b54b369b39f,
98'h0e10b3a1e160634093605b045,
98'h072c0c8f9838cddfabdc45b89,
98'h0b2a783b94d8881e67d9369bd,
98'h0410647560ef33440800c0168,
98'h0f30db4fa191f943e93fe5ee5,
98'h0b383b693074c65bac30b524e,
98'h0d05e6f34be6da830eeb40713,
98'h04248b7909116c8f663b305d9,
98'h0d33d46aa7b4891ca34d7e022,
98'h04060a61cc3e4737ad3a1761d,
98'h0a3c512b3896dcc1e41114666,
98'h0a18e68ff1f50c9db0b4cb7b4,
98'h013bf3da37fdd893af037ccb6,
98'h05193420727450faae4e731b7,
98'h0216e14c6dcecc22cde36146c,
98'h0a3d09e0ba01bf77cbf96b5bc,
98'h0e13a1866771e46fb10fb2561,
98'h01114e4e62a3432e0d61617d8,
98'h073924bdb25d2cece8ed245f1,
98'h0a063494cc782025ae65946aa,
98'h1534f85729de007a659f952ea,
98'h19a8699290cafc58cfc4be346,
98'h19beabe83d51ea68ea9cd97ad,
98'h0233f0d3a7e5d8af95c425944,
98'h051d6634faeff77a0a867260c,
98'h0c1db195fb60fa039003576bb,
98'h0424aa33097376deb1dfaae65,
98'h19a0b3c50155c21d636608447,
98'h002d4c071aa92b3786bd9d78a,
98'h070c0cffd80e78b5c6b59dcfa,
98'h043f9606bf0feb9647c6a16d6,
98'h183e7d91bcfc0476b0d3e0673,
98'h01139db6e72db47b154ea0821,
98'h042cbd78196a93f80a10548c7,
98'h0c3cc8cbb9aa28d78765d45c0,
98'h0d3f7960bede36c3f179bc68c,
98'h0505822acb2f830c13076c092,
98'h0f05ffa7cbf06651a40d414db,
98'h01301ee8a002f5eac6bd997e6,
98'h152a9d5a15377f0c284cc534d,
98'h0d01f34b43f57db32a9887199,
98'h0f05ab35cb71294ba43ddc3fa,
98'h002d97c71b3e2117a69db5206,
98'h181c4aa6f898b258e6daee37b,
98'h07215e0082bea238342d3f3ff,
98'h0407d2cacf82556cc278000e3,
98'h0f2ef5cd9de39fa604e28a0de,
98'h19b2ed6e25c474b14b44a55ce,
98'h1531423322812562cfddd887d,
98'h0b09640e52e7c23e0dec99e57,
98'h18055e654abcadde277c49931,
98'h0a279cd80f07591d48b08310e,
98'h0b1bd2ca778592fac64bbd7d5,
98'h1506c7a8cdb9c646b0a859714,
98'h0f16f9f5edccef0848b0237be,
98'h0c12bb0d654c01a4cf38fa3f8,
98'h0b1b95adf71dedc8ec57af2c8,
98'h0a0681424d07570fd08e60ddb,
98'h0b2893e691278d6c05c376148,
98'h0d1c9534f92b3f5007140854a,
98'h053b03c63638cf943191f5213,
98'h0a0fcf81dfb4291faedcf4d69,
98'h0c333aa0a6605a518a70fe286,
98'h001a0376f4383227aca4e53c8,
98'h182028fb00508925ed148d67a,
98'h0d0d4c10da92d000661c2c884,
98'h0f05df8b4b98ee0169e807045,
98'h001508fbea086932c6a7b3633,
98'h0024443508b64244aa875c8ba,
98'h0f1b8b96773ade382236a19e7,
98'h1832f70ea5e9c7c211959a73a,
98'h050173ebc2f802792f872fb42,
98'h0a37675c2ef919b9a1fe5d994,
98'h1803bdba475b054fee4c20457,
98'h0d0a1892d4276ddd07d7b0c29,
98'h0f1d7d6e7ae9cb03884c619bf,
98'h0c101757e029454c9281d21c7,
98'h0f224d25048735cf4b0e57291,
98'h199d9e7ffb038d99c4ea60bd1,
98'h013e69abbcc35eda55284b066,
98'h0c26ec0f8df731c52f8072217,
98'h19b97f7eb2c2bf3e468787753,
98'h0d14463d688a1b3fd31f0faf3,
98'h0f0927cbd26549040d67985f4,
98'h19be306cbc6ea2eb085b9c33f,
98'h19b0156f20067025558b34d5e,
98'h1986d033cdba72182e6da1651,
98'h0b16f1f66ddf2389e9d050930,
98'h0c358256ab0dd3874e3d85601,
98'h183bea9e37c2b60bcdd0d5777,
98'h0d299fca933c7469b3ffa82a7,
98'h0e05ed53cbdfb7736819850d1,
98'h012972b512f89560a6796931d,
98'h183895b4311dbd7a650882057,
98'h00025b6ac4b1ab7d325594cba,
98'h0535ca0c2ba11cc8812d01ba0,
98'h041f25707e4771404c35b9b52,
98'h022a0858942d91f81099a5ac2,
98'h0a298c7b1322679a8595e6942,
98'h0230634720d0da91e752fd056,
98'h053bf17037f2c6eda8c04f764,
98'h002b2f34166e3e0e0f4bae177,
98'h15183f64f046e009c5a65b508,
98'h0a3e5f2d3cb406d63157c7dba,
98'h1809009cd219ed3071bc9980d,
98'h0e0891ee5133eb43aa88bb735,
98'h1501a38ec36c531287cf1f4c8,
98'h0b27cee58f87669ec61b7da85,
98'h1982efde45e651d106abcd611,
98'h0c06f32f4dd9022167da506bd,
98'h0b38ab61317625fd2677fd543,
98'h0020ce98819b8df36f2bb4579,
98'h0b356f1caaca9997c06f17230,
98'h0f15f09f6be84a2e0d80022d1,
98'h0121ac45037b0511aebf8eb35,
98'h0a22256e846cffdb01272c55b,
98'h0f22e13f85ddc04be3a3c9526,
98'h0d2ea2e51d4309f345402862e,
98'h012ffea11ffe0397aa9c6b361,
98'h19ade58f9bf84e5ea84b808e3,
98'h0237fc2f2fd238b5ed698cfb9,
98'h0a1e3daafc4326f7cc828d394,
98'h0d2f9dde9f03bbd751985928a,
98'h0e000c23400a3a864b0cd66d7,
98'h198b68d3d6c90c9d438291aa6,
98'h0b3caf96b95945c46c151d5c4,
98'h0d1ac86475836f18d1257d56c,
98'h022b2151964bd459d0a78ddf4,
98'h0229631512c0fccac61dbd6ad,
98'h180f42515ea6e9e0053a97f7f,
98'h0f3b9f9ab73425a42dad8b0c5,
98'h0120d842818a9ae0d19bf14fb,
98'h042b59db16a1a10600aadcc8d,
98'h0b173a82ee5495d466b33eb84,
98'h0a19c7ea73b5cec12e5af415d,
98'h19a6af1e0d7c9c232f73e5aae,
98'h199b8f0df722881709c8d2d05,
98'h180c77d2d8e3eb27942f85c93,
98'h053408ba281660b86c3c18be9,
98'h0f368f0cad009529cb529a5ca,
98'h0024b795094e57c5cf0dc90d9,
98'h0f0414e9c83dca63225cc3d6b,
98'h0005ec734bf2f8d0a5d077d34,
98'h040b6c3656da11fc62fe39510,
98'h0f0d9b59db21ecda06b95f8cb,
98'h0c03076f463c730e2a8be20cf,
98'h1999607cf2f4fb53248fde9f6,
98'h0019e5c273e98da2132396f40,
98'h0b00b54241477b1c4d00dcd91,
98'h043cc00bb9b1a3b123120c17a,
98'h0424553f08ab33870f7b98ef3,
98'h0d34e5d929e092240333e2318,
98'h011fd3387fadad540dc55dff4,
98'h19bdca66bba8b9d3903360231,
98'h02325e2224bef3b4b559a10e8,
98'h199e41a2fcb1d889a9bc5475b,
98'h0a23b622877ac54a3594068b2,
98'h18026d28c4e4d1fe04679edb3,
98'h199a518e74853524c739cfc9b,
98'h0c035946c6bd68dab387e1acc,
98'h0f07b1e9cf5bbbc564b030886,
98'h183949f9b29ae7b86798db6bd,
98'h183fe8eabfebb81d92b50c6c8,
98'h0525b7ed8b78ba1fb60ae8420,
98'h15014d75c2af608e84279c835,
98'h0731fd80a3e7f58a05ec2b811,
98'h0a2160a002c223e8cac67cc2a,
98'h0b2fb3bf9f52d260e338e1223,
98'h0103e2aec7cd7a6dcaa0a1882,
98'h0d37bf672f4314fbc23457472,
98'h05311816221f26cdef1eb518b,
98'h07350de42a1466a569d40fb90,
98'h01103e7c6069e72a0c525d226,
98'h0f180254702b9e95085e89699,
98'h0e3b31b5366196140fd0e83a5,
98'h0c1f9283ff3bfaf5312731f24,
98'h041040c66093bb8cf2d6e35e4,
98'h021513efea1349de6928ff14d,
98'h0b1732e4ee4d8e04cb0a17739,
98'h1807b8c5cf5602596e59303a6,
98'h013e7c753cd0635ce9d76ec7d,
98'h0204bce249444d5f4f83b7f48,
98'h0025a40d0b4591e6c2d242906,
98'h153942d23290fed962dacd7cf,
98'h0a19d7717392c162f1f2906ae,
98'h151ae0d375c37e9fcf6b26351,
98'h0019b096735fac02f2b797dcc,
98'h0223ddd1878da17cccde57265,
98'h02252aa10a4e4f66c26c5fd39,
98'h02201e6b002e7228031cde81f,
98'h180ec6e85d968da06093a424c,
98'h19b7c1ec2faaea4b8d6955223,
98'h0c32e1eea5e63e301258ab0de,
98'h19946f51e8d59b806c864807a,
98'h182a386a9456af07709a82b49,
98'h0f2e52491c8e484ecb2039dc8,
98'h043c9c40b93895872aef26a5f,
98'h0f3dc82f3b926d306f5d4c71f,
98'h1508d985d1a76f8012b40d57e,
98'h003ebd10bd67b98d89ac12417,
98'h0506cb7f4d8554344f699da78,
98'h0722b8ab055978bfe4a307ece,
98'h0038a1a231703553231f0c5ac,
98'h0d3e9b6bbd31eb102c6a35bd5,
98'h0e105492e0b18ffeb29c219ef,
98'h07310b6e22088eb74bb079246,
98'h153e4b26bc998dc7ea4e66895,
98'h0f2e91809d2e58de1475f63ba,
98'h010e2f635c6695af0b173a97a,
98'h0c10661fe0f0de9e275d31449,
98'h0526f37c8dca4d264b40512f8,
98'h1532ee78a5dd6e0064bc5028b,
98'h043306d8260d090dcec4171e4,
98'h1520e96801dd16fd6a9003f97,
98'h19a5bb0a8b40aeb645bf80196,
98'h0c384c7bb0b2a47e29399a703,
98'h1802d8d9c5a404e10f3abc3e7,
98'h19a5d0ef8b93855be769b76eb,
98'h19bd6539bac774c0494e5592e,
98'h000430b14844a55fd521367e7,
98'h0732965025343af3221235844,
98'h041c135d781436426b19b450d,
98'h0a35f871abc7088bcf0c1267f,
98'h19b1ab41237968acad7f403f5,
98'h0413c323e79f140aef4ac4fb7,
98'h003d025a3a1315386aecb5cbb,
98'h041e5e1a7cb29a60ae9405e4a,
98'h0e19f754f3ee556d90343e1ec,
98'h020c163bd809cfefd08213309,
98'h042cea8d99ee0cc60685798ae,
98'h0b1a029bf41141886786bdd4e,
98'h18291b12121c61aaefcad1091,
98'h0a1919807224a56a8a915f2f4,
98'h1815b39feb5f2673ef0f6fbab,
98'h0d3a755db4e31c4890dd3684f,
98'h011e87a2fd38326b308764698,
98'h051fc9d9ff8de2434f95ae838,
98'h0b2d80389b2aaac9112b6b074,
98'h0f2508c88a226feb09960ac06,
98'h0739b92e334e3bb74651de2ce,
98'h0508372fd0510b41eea1fd395,
98'h18294e001289414e4556509c7,
98'h0c04724448e0c8b78aaca3d39,
98'h0212d6dc659ae09765394ebef,
98'h0125246a8a41fc2e49eb6ddcf,
98'h001b959ef70e108b42d9c8263,
98'h00066a38ccc019f5cdca698a8,
98'h051f52d4fe9e93136331a10ba,
98'h0f27a7728f7407d030ef797a1,
98'h153eeabbbdc8de07c7a6ebd0b,
98'h0b254c0d8a87ddedd4c1f230d,
98'h0d228a40052df432856b4a7ed,
98'h021ec92f7d8d17efc4941f9ca,
98'h052c9bff99242e4c0feaf847c,
98'h153db62bbb5635e767943292e,
98'h150a6546d4fdf3fdb424fb04c,
98'h0c0325884674cd552a8216512,
98'h0c3f53123ebf64e0249dfcb76,
98'h0d3029fa206d0a2a92bfadfc9,
98'h1837f70fafebf17c8b674d092,
98'h050e8b665d1f9fc87208fa230,
98'h19a1b49b8344e44c488b8acbb,
98'h0e0eabe1dd5b29ffe739a639f,
98'h02341dc3a801dab7cada75787,
98'h181f9cb17f35fe112a8d7e1ed,
98'h05090044523c2e1835d566b0a,
98'h0e166349ecc16bae45d14b972,
98'h0a10228a60764cb62eb5f3be0,
98'h19a96e5092d76df86aa19bd02,
98'h021bb0b2f75802cb6b2037124,
98'h04353a9aaa73cc7f2e5cecdf9,
98'h0f32598b24a8b3800baa41c67,
98'h0a2f282c9e79ac442cf6c342c,
98'h0d041b90c80081eeca2a351c3,
98'h0b1b7f3c76f690b92541275fe,
98'h0e0ec1ef5d996a1e708483fd6,
98'h0c0ba52dd763ccbe8aea0b037,
98'h152f11851e194a0968dbdc7b1,
98'h18198196f31763a56cd216e3a,
98'h040ba5de575dda9872cc394f1,
98'h1805133b4a055a2ec6da601db,
98'h00367e382cc398a448829b5a8,
98'h0e093511d262778b0b3e85b71,
98'h19923a7fe4509df5e81aeb273,
98'h152c933d9929765c0f78b61d7,
98'h19b80852301c6a466b9582666,
98'h1503d01547b3a5b2b2751ca62,
98'h0d0b3ffc567d9c3f272ddd720,
98'h1809d91d5385fa0fc8e2370ee,
98'h0217b17aef769a78aae3f4cb4,
98'h02236c0a06e38e640c6392fce,
98'h1987a17b4f4a2c7c4241be9b8,
98'h1992cbc165a695108a34737de,
98'h152e765a1cd103c26fce58347,
98'h0510a5576150b8e76c7fde872,
98'h07151524ea1934b4e998578fb,
98'h19af25119e73ee27ac4b92767,
98'h0224ee9809c89fac4e08c4ce5,
98'h0f1c3b65f844b38442fb63911,
98'h0c3ebc213d6b49f111d83bba8,
98'h198811f75016c31cf26a81848,
98'h0039ecdd33c6a6bd4a67b5451,
98'h0f24b09c09753382ad0024e69,
98'h0a39c298b3bad039a6267907b,
98'h0223d25987b708b72f7d24b49,
98'h04351ed0aa2ab07e8276b6c43,
98'h0a07ea63cfe1352a8b97f3d3c,
98'h0a3dffb2bbd41a95e67a47e39,
98'h0f0d5920da970abf718486922,
98'h0105ad1b4b70d3772a6918f81,
98'h0f20d124018a1bc4c31da024a,
98'h020a9597d5298b0d042abb3a3,
98'h1507ec344fca8bfd45cd08293,
98'h150cdb64d993c53069349e0c6,
98'h0010f04561c8d198cba828255,
98'h1816916f6d23b2a8887670778,
98'h180ec47cdd89e638d14e9105f,
98'h0214a854696afa300d662aad6,
98'h0216162f6c3ee7ee2adfe8a11,
98'h022d8b611b2d71700b953f876,
98'h19a0ade181612a3a0756bf344,
98'h04326d9324c4c600c6c07606e,
98'h182bf44997e3b70d8a3dcce4f,
98'h0f38469630bc166b2c03ead5c,
98'h1517a74bef7b3fc92ffd17405,
98'h01157fc8eafc7b28b124b9c54,
98'h0739befd336d7e3e8b047ebc6,
98'h0d31513622937fa1eea9cf4ee,
98'h0c0c82a2d90905ae4bf134360,
98'h1981ce9cc38c8b30494562144,
98'h0a0bcdb1579683c9e74396734,
98'h0c05a468cb463a1c4868945ed,
98'h010684ce4d0471b145d2f7a14,
98'h19b684b7ad1ca69fe382bd9fe,
98'h01193ace727e34f631b4cad5e,
98'h0f21445602b1a1e2ace5dbf12,
98'h043705b62e0fb099c474b98e3,
98'h0000a7c1414bdcfecc91ad93f,
98'h0d1583bbeb26460c005321300,
98'h1527e0260ff601fcae0ef271f,
98'h020110434230462fa9477888b,
98'h0f39b861b376bcd5a10c559cc,
98'h070e28e25c4bd254d0ac1d4dd,
98'h18197200f2eab47208d67ecdc,
98'h0a0d025d5a262d3b92c1099cb,
98'h0d325240a4b973ac290ccbe63,
98'h0f144da9689c7c166c7af17b3,
98'h0f22df0e058e424bcdec326ff,
98'h0c282ceb905ef785652c48567,
98'h1808cc06d1adee0a8721c91c4,
98'h0132587924878c99ca6dae845,
98'h0f1a9776f5328391296e7944b,
98'h073073d6a0c4edd4d11346c20,
98'h002bd75b17a5f77889fd586ad,
98'h052d92b99b2b142705f473b4e,
98'h072936619264bf4a081629b82,
98'h0a0bee06d7ea2ff206637d6ae,
98'h0c0920e6d2615a7e887d877e3,
98'h0513c8d3679d0a06679a9ed95,
98'h151e21f7fc51cb7eeb2c34b67,
98'h022c8563190fd4a4d45bfb5db,
98'h0d27f0508fc000a446cf1681f,
98'h0114ea2d69d06c7f6739fc3d3,
98'h0c302b6020662d370ab955ab3,
98'h181f96d4ff0909b5cb259625c,
98'h052fc8419fb01271b5ca2822a,
98'h0528a92f915660d9e937f6acd,
98'h0c2a2ec3146a387b859fc2826,
98'h02299243133a33ec282519cfa,
98'h001b0661f618176ee558f18bd,
98'h00001b43c03b535e2d8cc7743,
98'h1803b349475a3053e00edba88,
98'h182d9a961b340f1027d778e75,
98'h0c158357eb3d1623acd86a699,
98'h010358cfc68017544dd4a65ee,
98'h19a58b1a0b3a66c721e0dc090,
98'h0a2125b5826acdea0937fc785,
98'h0c0732cd4e64b4180322fce7e,
98'h199b1d3d762f0703869af9b95,
98'h071a735df4e75cde93f289103,
98'h050b9c8a57093a41cf00740f1,
98'h150ac36955b355d4a70535b30,
98'h0e0666f2cccd23b54aaf864f8,
98'h0c2bb43c1761e2a206b4e2aa0,
98'h0111fafbe3dfd4df68e365b78,
98'h0b103ed3e0463ee0c93c73f6d,
98'h19bc1759382735b08ad59f6d2,
98'h19a9c0dd139737197478d3426,
98'h0e0e6ff1dceff58a8b503dfda,
98'h022ba9b51749b1c4cabf995f1,
98'h001892d8f13aec3da65d56de7,
98'h1520d76881a5284b8c54dfc5a,
98'h19b3fd5427d2eb0be5b17fed0,
98'h180fa3b55f4b10085061ba180,
98'h0c1760d8eefbfda4add6acef6,
98'h0d39a107335a33426ec4d79f6,
98'h19be180bbc3d1b2a3024f5126,
98'h0b34077c2806fa33d57ecccd7,
98'h0418cbc1f1b5472d2ccec06bf,
98'h0405d1e0cbb1a404ad7384bbc,
98'h0d2c4800189d22aee3eddd796,
98'h0c288ab191336fcea9725aabc,
98'h0d3380fb2705ed1fc756fea01,
98'h0438c91cb18bb59acd0e5b86b,
98'h0c09c818d396f560ed711fadd,
98'h02135dfe6685ef61c7e82f5e7,
98'h151230ede47a7ac3aa2653580,
98'h0e0c30e3d861b20c8e632aec6,
98'h0d01263ec25afe08e99b78bc1,
98'h199bcd0977b5967423d70911f,
98'h199d2f00fa420261545458df6,
98'h00109e5d6136126234f7cc588,
98'h19bbe35937d93e6ee851ac2fe,
98'h1500de7b41b9418eb46548720,
98'h0e30119ca03f3d4125ae88028,
98'h002a31b114409ea34b9bd3b77,
98'h0c0e13505c106f59e51ab4151,
98'h051bf3fc77c1ac38ca07a0aa9,
98'h071b522976b5abaa2f37680d4,
98'h0b39360832568dd86f743f74e,
98'h072dfd0c1bf920932f63f0f82,
98'h150f6a335eef90fa88c9c767d,
98'h19b1ed0ea3d2b4e56cffbecb7,
98'h022ec18a1d8ea6094f61287d0,
98'h19b7ba752f4cd8e247ef59e4d,
98'h0a2138c98245c95c524124d5d,
98'h19a301b48612c73a6319c0897,
98'h0f0d555edaa15c3d87ed723bc,
98'h073cd872b9a9360e8a6bac671,
98'h0c019266c3176de5f03983a04,
98'h001f7283fec277f0c3c640133,
98'h00157dae6ac4f47dcfb87a9d2,
98'h051ff6ecffcf0ce14ab69c8b0,
98'h19bd84b23b31f61eb13bc0f38,
98'h010b84e3571ba351753bdeb43,
98'h071e71a07cc5a1d1c609ca0d3,
98'h023c68cbb8fd892130f904dc8,
98'h011d9854fb03588fcece7c7b3,
98'h0a3c813bb93e8ca32f083c392,
98'h001ab35cf559a641f0dec377b,
98'h0e19d3f7f3a94d970d5d1667b,
98'h003070f5a0fc2ac03070c863b,
98'h010252f4c486fe2f484b26ed7,
98'h0a08b00c517172d5216254490,
98'h022bd157978f940b46de88b86,
98'h01016d3dc2edc138866ed958b,
98'h0e3d2876ba7d693ca0fbcb9d9,
98'h070f5fd6de83c794522ea46cd,
98'h0c1d8cd57b254d448964c9dac,
98'h153b46d436a44f8091d0b6867,
98'h0e3f13293e24061392f7e5952,
98'h0406e5e3cdd5d3877318c64f2,
98'h0429655712e2410b84772e5ad,
98'h0a36b261ad7d0820a5c2e998a,
98'h0739a774335ff3fcedeceea09,
98'h152d305b1a7f54b62ea666dc4,
98'h003c8cc5b9282e288beb21445,
98'h0e34ff8da9f83ca02e592ebb8,
98'h07379cc0af3e593fae0b4f0b7,
98'h000698664d2ab8288d9d7d801,
98'h0526a8090d45ea63434c5423b,
98'h0b06b900cd477d87c49b249b1,
98'h0c226d7504d5832466138da22,
98'h0b2a822b151139e6e43dfc266,
98'h15156f09ead68283e80eef048,
98'h0d1e44627c97ba5eeffafc637,
98'h0113f6fb67c205f2d26d7fb05,
98'h183bfcd337f304f8aa357f3b8,
98'h0f1c4caef8bc5a52340bc072f,
98'h0f0e825add1761adf1f629c04,
98'h19b419b9283fdcf2ab0979023,
98'h0e0e62865ccb5366d07cfdaaf,
98'h0c07fee04ff84c95aab66d7b4,
98'h0e356e922af880fc270012dd8,
98'h0a225918049f8a6cee4b7be39,
98'h0035f86babc08e3843b078e14,
98'h153e3686bc5ccb17eafda1a8f,
98'h1812bfafe56ee4d29466c067a,
98'h072b7b8016d737a86f6069209,
98'h0e048eabc9106d756780acca2,
98'h0129378a125cfe9f65c53f085,
98'h050a875cd52a38b884e18d8a6,
98'h0f0b2a58d66fd4ed068d30055,
98'h0d32206f24781826295ebfd17,
98'h0b2f78d21ef7e6f42c6a8e255,
98'h0513d240678c2736ca89d7f19,
98'h1539920a330e3984cb27fe5dc,
98'h183173dca2d844537211f2e3b,
98'h0d374446aebf7adf2ec26e0c0,
98'h04134802669a79d46efdafc97,
98'h0a0501fc4a1843b56aab7075b,
98'h0b30ba1d21555703e507516c7,
98'h023656d02cbbc827ab2184484,
98'h0f21cb4b03ad39198bbc87bdf,
98'h01378c972f35f8c7a4b3c1192,
98'h0c062f58cc73843fac1b6157b,
98'h150d80565b2a1396061e6ce62,
98'h0b3f19c2be18cc8eec0de4fb1,
98'h0508a742d16ea5041255f9946,
98'h1508bab6d16eef0f859dd311b,
98'h023043c12097f8f2e99dea719,
98'h15306c1120d41abbe8b20f2d0,
98'h0e1aca6775a1fbb20d8121b34,
98'h0a148e5f690fc97bd0ef31865,
98'h051876f970da8b04ecc915f6c,
98'h0d0b15de561aa9286d7cc07f9,
98'h0005116c4a1d371a68c96fc1b,
98'h073bc77ab7ba748b22889221b,
98'h1985e2e5cbe173940fbd8f017,
98'h182b25d2164abc5cc959d59e7,
98'h0128daba118c3883cb9d788bb,
98'h07230e31063ba04624ad44cf7,
98'h0d09e36ed3e613698357ab9dd,
98'h0c160594ec3f77e0a83bfdb61,
98'h0c1367b8e6c6a8374e155f5d6,
98'h020a35aa54506bb56cb683fc0,
98'h011f077cfe36a24ca596a857f,
98'h040919ce5226fe3c8fd56a726,
98'h19ab7cd016f9157c258c0602b,
98'h0200dc0e41aa84e00c2924931,
98'h180cb0f7d95d4f05e0ead83b9,
98'h00346226a8d490f8ec5a7fff7,
98'h0a2b0168162a169a8a423cc7e,
98'h0b070a84ce3048cea8154600a,
98'h0c16b4c76d635f5c864dd4d4e,
98'h0f211945020eb09bce5e8508f,
98'h0e249fe9091b68dbe44bf2783,
98'h1999d535f3b8e388a5d002314,
98'h0b38fad331f05018b354ae2fa,
98'h000454d348993caf6f4a52baf,
98'h0f1565baeac71085c2276460b,
98'h022bfb4997c47016ce771d902,
98'h152f1e041e04f503467c1ad81,
98'h0f3da577bb7b93b9accd04c1d,
98'h0202634544f878e1b2ae4e4c5,
98'h0d0a86e8d5301880a1beb709c,
98'h0b080c41d01298e3688ea7da6,
98'h0201b6dac342b344c6c6a9495,
98'h04224bf004819437c1511a87e,
98'h042d6d3a1ae635ce0228f809f,
98'h0005a6744b6e1d8087c4e8c20,
98'h0430efa4a1ff57d6a2dcf0fd3,
98'h19931623e60bfbcf498c11ded,
98'h15342e66a84a7007cfe7c47cc,
98'h19886083d0df1ba46f5fa79b9,
98'h181a117d74001cf94a99df0a1,
98'h0b1b9b48f7060ff0d3068b9da,
98'h070e7595dce1de3490886ace6,
98'h0706e157cdcb031548fc14f29,
98'h0128d90c91879d32c534791b4,
98'h053937c5b26c17e384ac1d8fd,
98'h0710b8ef6177265d2de953ea4,
98'h0111a2d8637c3a9c2a21f7d32,
98'h02009dfac13e920ca923775d2,
98'h05396b0432ed61f080cfcc01e,
98'h0734d99ba9ba9d89ae09b33d2,
98'h052291ed850540014c3bddc95,
98'h0e02f2efc5e1f40d8289f47bb,
98'h011f776afeed635f04f939bf5,
98'h0506c3c34d9e67c2700336b27,
98'h1838ae80317fc80ba4a94ae17,
98'h0d02459344ad1abf126e1da2f,
98'h0a1602626c20d877046bd8149,
98'h0a3d0e8d3a2e980e0d8db6b65,
98'h19bfab773f67de83911ae9a6c,
98'h0a207e8d80ffdca7b649e27ea,
98'h002cb4529946e48142c816cd5,
98'h073d9c223b255075865ce634f,
98'h0d038ebac7130631f098bb25e,
98'h0f19a1877340af50c505a53b3,
98'h1521d8a383be31c5309694360,
98'h0c0e39a9dc7ae2012638029a3,
98'h15305133208358dd4a2246eac,
98'h043a6d26b4fac740ad6cea841,
98'h0c37fdbdaff6118aae4d4d19d,
98'h18313f4ba271ecb8af0b83d21,
98'h041d7ec87ad6a74eeea8cb011,
98'h1502fb15c5f838012fbd0985d,
98'h0e1795086f3b9c1a26beccc5c,
98'h0d2e30309c5f7fa3ef54cc48a,
98'h1525d6620b91994dea636bf52,
98'h18355ffb2a981419682ddbec0,
98'h073c92ebb922d0bb10b35d052,
98'h0f065a80ccaf38ca1017d8e9a,
98'h0a0ae9e955c6cda2c6ed64d2b,
98'h0b104b7f60a08d1087f46de30,
98'h18300ecfa00bb5b64aec3623f,
98'h021577636ae365348e0ef1217,
98'h0e24be448959fa15eb3e3725f,
98'h0035a84a2b4d137045dfae16a,
98'h020de31cdbc37852cae0aeee9,
98'h0c1e4b00fc9120eb677456dbe,
98'h0b1d6b5cfadf0b6e722bdafb1,
98'h0e3d3c03ba5876bf717f1db2d,
98'h02164d3a6c818cd8d2256cb0c,
98'h0f034480c69876f56ba5f684c,
98'h0f38bc19b15545746566eedd9,
98'h0d33475426830586502380638,
98'h050b8d90d700ce914ced93369,
98'h012b1e0b1618815ae70317088,
98'h0527ce638fbe62f025d0e7d98,
98'h010325e34654ad4ce5398c54f,
98'h071b8787f7349fc2a1d5f4cc1,
98'h01117cc8e2df89246f9409d2a,
98'h19a8b3221151b5a9e8fc417b5,
98'h000dee595bdb1a9b6abe9a330,
98'h18156187eada09b666fa423d3,
98'h010390e147172659f0bbdacf9,
98'h19b20e3d240b46694206adced,
98'h002d125d9a23d8f90f6f55299,
98'h072b24f81664dcb386943ad5a,
98'h1988b57c516c60028764006ae,
98'h052ab69d1556f4f6eabd455fb,
98'h0a20fe9901f272ef26a06ae50,
98'h013f5e41be88d002c304dc621,
98'h0b3710c22e33cc272ff20b911,
98'h152d56299a9798196e5ab73a5,
98'h182bbab317729204abf13b90c,
98'h0f3ebccbbd5ea1ebebe7932df,
98'h0e3433daa849afcfd32757ade,
98'h0f1809cb700a1d9a4d9f78ea9,
98'h199789546f261ec20fc889d96,
98'h1505b2fe4b6537b6122f6a059,
98'h0d21baed836e1f04081abaad1,
98'h012801699004aa40c423f67c6,
98'h0a298824130f60af444b2aea9,
98'h0a121642641ebdaae74e3a34d,
98'h0535ed23abdd1ccc6b8c34fb5,
98'h05211fec8211b9d4ec44c27c0,
98'h00004fca40971e5461ccb6706,
98'h1800befe4149c710c025db87b,
98'h0a005ca4c0a2bb2f8652a183c,
98'h19819b3c43273f1e82a8c5f51,
98'h071e93effd2ebd38872a3696b,
98'h0f17289bee766e303113544a1,
98'h0a1a8698752b3b370f6365b30,
98'h01019c40c339c3e62fd17073d,
98'h0421c33b83ae61e5010ed809c,
98'h0419118172377451a1f409482,
98'h0b047326c8cf2ceacd942174c,
98'h0b1edee27dab88f384f4e8046,
98'h0c24a756096f0fe1123299f57,
98'h0e2a1b17942f61bd0564edcdc,
98'h0a2d55779a9b8f51e8965f352,
98'h153452082897a60f693239326,
98'h198e04e7dc20c9b50f72fe05e,
98'h003b69c736f9a5ba2d6bb3a73,
98'h00282bb31055f0746dcd43e05,
98'h0c1db79afb792a00241f8709e,
98'h0a0b3b97d65cb0e8f1e5b866c,
98'h180544f74aafb6910819fb203,
98'h0b0c5f01d8bc8d5aa8ad3ee21,
98'h052744820eae3a8e88f23b172,
98'h0436e60eadf3260424f55fc42,
98'h150cb710594a3189cc8a8304b,
98'h0f02638b44c2720d4b95ba268,
98'h0b0940a6d297348364f135662,
98'h19ab79f416f5e88f27681d4a9,
98'h18352d79aa5dfaec6c2858a0d,
98'h0c3c58773887999350a4ca198,
98'h19afa6ef1f51cba57130fc829,
98'h0701e7f0c3fe37122e405ca52,
98'h0a1e189c7c355e0022c007c0c,
98'h0d1aa7ee754d0df55194dda72,
98'h020dc5455b902abd7099ed78e,
98'h0e3c3babb86eef1487677c00b,
98'h0b0c8bdf59052d0dd1aacab00,
98'h0f3ca717b965083a89046e3b4,
98'h073ddc8fbb8c139352286bd48,
98'h0f1c3bcdf872ad1f30b27c08b,
98'h0f20ddab01bde15db1e3ba3b4,
98'h053d361bba5f106be437afc23,
98'h0c2cc0b69995feee6fe711a1e,
98'h0e2609fe8c35ecb92970afe94,
98'h01184767f0b8bb36a696fdadf,
98'h021b6022f6f01d90ac7440a7a,
98'h199178a2e2c03c97ce42df6ce,
98'h040ec2e5dd9d286b6f146d4ea,
98'h0c1a857d7500e1e1c86afad45,
98'h198efb54ddd6b5b1f046d9d7c,
98'h0730de3ba1a613568dd96c41b,
98'h05171e2c6e36f9bcaa35bc648,
98'h0a13775366f883a6acd385fa4,
98'h0e0948d952bb0dd62c42febe8,
98'h0b2d3e691a4ee0f3483115abe,
98'h0e120e79642a3936095f07d71,
98'h0f18bf527159f5cd6c8f11ebd,
98'h0c2194d8830b2a06501cad47f,
98'h0121f91303ed3a3583cb2fb7b,
98'h0b176174eee01e5f0143ccd22,
98'h011b62e1f6d4d49dee7ddff4f,
98'h022dd67a9b92fd4a6dfc0ddff,
98'h0f0b2122567a0ae5a77034f14,
98'h05225fc704aa5fc009614b020,
98'h07256a6a0ac7235fc2732fe1c,
98'h0c074fe74e9089aa647b23727,
98'h07391c7e322bb5cb86a5f6647,
98'h051c6d1878e552e08e5934926,
98'h1523815307126c5bef806ffe3,
98'h0d3b2e46b644002dc70d7b6bc,
98'h0110440e608934afd0dfcb9d1,
98'h0f13a81067560c4968665e2f8,
98'h0b3a9605350ce0d94d9a6d167,
98'h0b2729c10e7be0dcb011ddb79,
98'h001483bbe91938596668c2a77,
98'h0c1d8a56fb047f814a4b6f055,
98'h0e2979e792ce792051c882760,
98'h0d02257e445d1abfe83dfcc1f,
98'h1980fa6dc1ed48900457d00f9,
98'h0d2588940b119f1166db90bf7,
98'h0b368162ad1a1479660dc9e96,
98'h0f10cfa5e1a72bde8e1425770,
98'h182b9a0c1708e41d4c2dfee11,
98'h0227b2700f497c80cbcd1f8a5,
98'h0b2923df1262992c045c4bbc3,
98'h01064160ccb441412762ef42c,
98'h0534c77fa9a4a0c7836ea0a88,
98'h0b1752936eb168582bb65a11c,
98'h040f9bc3df2c14808e722ebae,
98'h04109ed5e13556ef28ceec111,
98'h0202fab045cd4b5849517d714,
98'h0e318ea4a312121f61f411822,
98'h0a108679e108dabf4c50e8310,
98'h0411b72de36a57f10ac6584e4,
98'h050a5e85549f0796e9df03c7b,
98'h0f3c074d383da85e266a59871,
98'h0d088467d132a72f31de6bead,
98'h0e03a490c7563e4f678ecae5c,
98'h152070e680dc704a655678b81,
98'h022f78349ed1f89ce57f384c4,
98'h1833d8f6a7bfbc1928405c346,
98'h02096c2652ef33108ffce543f,
98'h199ba2bd7761b73c053e27cdb,
98'h0c0e58025cb68f63343f567e5,
98'h0e240a8e883402c4aa3139d96,
98'h042b9e16170aae3dc5960354d,
98'h013ef7f0bdf3c533a6cd9314f,
98'h0727785f0ed6d8396fccaf491,
98'h00018297432e2b79857f94262,
98'h1800f589c1c596dec0cbeb843,
98'h0431a768a36b59f88671a31a2,
98'h0c04a5f2c9583da769e740584,
98'h01192d78f270cd81255738e69,
98'h1982f8a745e862fb8ce27ebe8,
98'h1802bb0d457c2c53a7dad6e8b,
98'h0b054864ca8c4934c75fb9d84,
98'h07361a9aac078721c56464666,
98'h0a0e9897dd07379c4ccf686f1,
98'h0b38afc6b1580a0c69c5740d0,
98'h0d25025d8a1ec36a6f242e74c,
98'h0b071c65ce081da445d0f1720,
98'h1990d183619e08c86643ce828,
98'h152d157c9a2df7ea8ecbb692f,
98'h19ae51851cbfd3cf2bd6c359c,
98'h0f10684160ef9d508d9b89551,
98'h071f4a917ea8b9880c0001647,
98'h0b342f17a84551b7517201065,
98'h0e192e83f24a20ec4cde6033b,
98'h0b293695925b796ef018d3dc0,
98'h183cf5e9b9f73be427612c012,
98'h1810927fe134ea39348d0c737,
98'h0d15ad00eb64f0488e515f2e4,
98'h010562cacadeac46ee1ea7525,
98'h0c0ab0b5557db0e3a2f903c47,
98'h0532c89c25b62b38a86218664,
98'h19829ba4c522466d0aba3cf53,
98'h198b0b48d632d72027a938847,
98'h19a3e31b87e0888e8bef789a4,
98'h1504ed5549d4357e68611aea8,
98'h0d102417605906e167b648b4f,
98'h1834317728456243cb5a4abe3,
98'h152720448e7ca1edb01e64eeb,
98'h02024f9344b700d128e8f08c9,
98'h150e6b00dcfb142d21ae54192,
98'h0f3c59beb8a09cf88c825fcb8,
98'h052ac65895ab6b0891f73dadc,
98'h041b113e760a7bfa46b58c584,
98'h0e28300910676fd90e89634e2,
98'h151a2b86f470dd8727a3e7f88,
98'h0b1d9e7f7b0300e75262c2438,
98'h0b23c73d8781acc1518827d9a,
98'h01096dd7d2f85a6c24a95cffb,
98'h18051137ca25a138050072110,
98'h00137ce066d24f91688aac9bf,
98'h0d111979e235cfed29b9731c7,
98'h19b1fa15a3cd736fcbd1ba59c,
98'h0c06d8394daeac520f5fdb615,
98'h043de0a43bd9320f666d6122d,
98'h0d3f62dabee179479005c4ace,
98'h0434256a2851d96a730837088,
98'h199950f3f2952a1e6b217fb52,
98'h021093f3613c9269330b9ec49,
98'h0b0651484cb7b397a8d349972,
98'h151f5b7d7ebe49e525ef81380,
98'h0d0feecedff0cce434f76958a,
98'h0b124bf4e4b689a6ab402eecc,
98'h199885aaf11720a56bf23566e,
98'h0516c2f76d97416772abe9941,
98'h0f0d68325af8edebacab8117b,
98'h0f1948d172827fd04a8195878,
98'h012f33ea1e591938f066f2286,
98'h1993dd7fe7a71b7987e21348c,
98'h180556874ab1ad7d304ebe3e5,
98'h0e33f5b027c54bed48adc1012,
98'h0b01c2ee43bccd19ad7e50675,
98'h051527bf6a7432a323afa4020,
98'h1509d63453b512e02be25698a,
98'h0d3d88b9bb315405aa2fba452,
98'h0c096c9ed2ee6310921bb72fd,
98'h0a38b95d3173006d27bdf3ebd,
98'h002526a28a582c5d6eeaee729,
98'h001ea3167d66ad22029f54c00,
98'h0010dde461aa18e58f61540e1,
98'h0202e50245f43d5e286ebdb27,
98'h0d3f4a393eac2f3b81fdc8982,
98'h0a39f0edb3cf3b4ad2fade5d2,
98'h010fd6a6dfbb63602f824b0e1,
98'h0010d855e18f00ffc832ce81c,
98'h0b0fa660df5b97c3e867f6556,
98'h0704c967c9b6d186aa9acf893,
98'h0e12c9cde5980e48642ee6bba,
98'h18373c002e46e1d84ceab6059,
98'h199aa3817563493d919f87761,
98'h010bceacd79f51de73bf7b2fb,
98'h012e7d411cd75c66662ac822d,
98'h010cd3a9d9ae157107817669e,
98'h043b4d0236a7adf186aeba46b,
98'h0a238de40710cd59eeb8bebce,
98'h0b3fa9e9bf452781c44d16cf8,
98'h0c211df90203905152a1345ad,
98'h0b38f14c31e5d72703892b929,
98'h0f051f364a25a4010f47b21cc,
98'h02369baead110063664ab0cdd,
98'h021ef4987dcd2601cbd1e7048,
98'h0e28c1c691809d26cffb06a68,
98'h0d16c5cb6d92a4dc67ea57bb5,
98'h042ed1789d994ed26eaa5aa9f,
98'h041b2c2df66da90988720812c,
98'h151b72da76e9bf378ea2354dd,
98'h0d208fcb012b2df293014c847,
98'h01129d2fe51271976392ef6f6,
98'h198f3461de770af1298943b1d,
98'h0d16dbee6da703a28e018fd4c,
98'h052cf65d99e14c4d0eaf77e43,
98'h0c0ac3bb5589de7a47c390aaa,
98'h013fb7dcbf787c40a865288d6,
98'h051b976b773357af302e0d075,
98'h0a157dab6ac1dbf3cf13bbc6a,
98'h0b3a1d0334054242cd35d667c,
98'h000f3c465e488c7fcfcfd7d17,
98'h0e36a2b8ad7befa52795f2318,
98'h023b54db36aca7ed8eeca4977,
98'h150533f04a7da0b8ae39ff322,
98'h19bcc246b98b4a36c7e0b52a4,
98'h051efe3f7df966cdb4d2031f5,
98'h19abf61597c88a4350c619434,
98'h0725e66a0bf674a4ac5d20163,
98'h010e6585dcf462ed24c716c3b,
98'h041f4d667ea4df6f0780b21cc,
98'h0131c68323b38bfcb0b10b355,
98'h070b0558d630cfce2939549ff,
98'h0427fcab8fc5432bc74ef549c,
98'h0b0b769656c922d2c4fb4ff5d,
98'h0d10b64be16f05220875265a4,
98'h1983f4a3c7fa7afdab9feedb7,
98'h040db9605b473679c85f9be86,
98'h0f024336c4afc14007d53bf68,
98'h022ee0969dc7bcbb44ec811db,
98'h05384b33b09915fb67fda7547,
98'h0c12c84be581875fcd74584bc,
98'h0e3affb035ea31ff0c6513eae,
98'h0a292b8c927a08cfb1094c6bc,
98'h182b72f016d1378de728cd171,
98'h0e33f115a7eb9f650bbf2a9f8,
98'h199f1b6a7e36f3582d87e41ea,
98'h0513e85567d1ee6875f583b0a,
98'h0c0c48c1d8898d7ecb3975af7,
98'h051e3666fc5b2712e92575902,
98'h012fc8cc9f82aa92d05e575e7,
98'h19a773180ec7418cc82c9cd7d,
98'h0010bc906149fc954a1bad293,
98'h0a2175e682ee25ef8856ae496,
98'h0d379d40af0543f74343e6f58,
98'h1518d2fe7195c544ef0f384df,
98'h151d71437ad6c09971aba610d,
98'h000f083cde312284b3fd0c773,
98'h0208312cd07b12cd27900ab06,
98'h0d1e5a2f7c914b9864a0d0fe8,
98'h0d395cc2b2a78c53126be971f,
98'h1804611248c142594ff83a456,
98'h0503bffa4779f15ca83168dae,
98'h012045d280b5d58fa31f6c55c,
98'h020d67f75afaa98aa07586d89,
98'h1821af0e036a69f5874204608,
98'h1832c80fa5a260ee06e30640e,
98'h0c155e116ab3b3332f754a3f6,
98'h07300ec8a00419084db244512,
98'h052c7bd898c15ce1c9cd09f43,
98'h1525aad60b6ca9c9877b762e9,
98'h070b96125737a38a28249527e,
98'h013d001eba38b293a790ce672,
98'h0f1e4c1a7cb9dda5aedd6cac9,
98'h0e224cb58491fb36f2f60a700,
98'h151cabfdf96ef49c84ad11fb2,
98'h0538bde1317544f4b3a2e8269,
98'h071f3f7a7e78cdc92dab80b57,
98'h041db515fb518b7df1660350e,
98'h0f0ec8fc5d87a3734fdbd024f,
98'h0c003cf8c041b5f34b259b1be,
98'h0f2cb0a119624dd483107cbb0,
98'h0701ae5ec351b7e66a23bf9d6,
98'h0c212135826c7c158294d9915};

endmodule
