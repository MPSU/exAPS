`timescale 1 ps / 1 ps

(* STRUCTURAL_NETLIST = "yes" *)
module instr_mem
   (addr,
    read_data);
  input [31:0]addr;
  output [31:0]read_data;

  wire [31:0]addr;
  wire [31:0]read_data;
  wire \read_data[0]_INST_0_i_1_n_0 ;
  wire \read_data[0]_INST_0_i_2_n_0 ;
  wire \read_data[0]_INST_0_i_3_n_0 ;
  wire \read_data[0]_INST_0_i_4_n_0 ;
  wire \read_data[0]_INST_0_i_5_n_0 ;
  wire \read_data[0]_INST_0_i_6_n_0 ;
  wire \read_data[0]_INST_0_i_7_n_0 ;
  wire \read_data[0]_INST_0_i_8_n_0 ;
  wire \read_data[0]_INST_0_i_9_n_0 ;
  wire \read_data[10]_INST_0_i_1_n_0 ;
  wire \read_data[10]_INST_0_i_2_n_0 ;
  wire \read_data[10]_INST_0_i_3_n_0 ;
  wire \read_data[10]_INST_0_i_4_n_0 ;
  wire \read_data[10]_INST_0_i_5_n_0 ;
  wire \read_data[10]_INST_0_i_6_n_0 ;
  wire \read_data[10]_INST_0_i_7_n_0 ;
  wire \read_data[10]_INST_0_i_8_n_0 ;
  wire \read_data[11]_INST_0_i_10_n_0 ;
  wire \read_data[11]_INST_0_i_11_n_0 ;
  wire \read_data[11]_INST_0_i_12_n_0 ;
  wire \read_data[11]_INST_0_i_13_n_0 ;
  wire \read_data[11]_INST_0_i_1_n_0 ;
  wire \read_data[11]_INST_0_i_2_n_0 ;
  wire \read_data[11]_INST_0_i_3_n_0 ;
  wire \read_data[11]_INST_0_i_4_n_0 ;
  wire \read_data[11]_INST_0_i_5_n_0 ;
  wire \read_data[11]_INST_0_i_6_n_0 ;
  wire \read_data[11]_INST_0_i_7_n_0 ;
  wire \read_data[11]_INST_0_i_8_n_0 ;
  wire \read_data[11]_INST_0_i_9_n_0 ;
  wire \read_data[12]_INST_0_i_10_n_0 ;
  wire \read_data[12]_INST_0_i_11_n_0 ;
  wire \read_data[12]_INST_0_i_1_n_0 ;
  wire \read_data[12]_INST_0_i_2_n_0 ;
  wire \read_data[12]_INST_0_i_3_n_0 ;
  wire \read_data[12]_INST_0_i_4_n_0 ;
  wire \read_data[12]_INST_0_i_5_n_0 ;
  wire \read_data[12]_INST_0_i_6_n_0 ;
  wire \read_data[12]_INST_0_i_7_n_0 ;
  wire \read_data[12]_INST_0_i_8_n_0 ;
  wire \read_data[12]_INST_0_i_9_n_0 ;
  wire \read_data[13]_INST_0_i_10_n_0 ;
  wire \read_data[13]_INST_0_i_11_n_0 ;
  wire \read_data[13]_INST_0_i_12_n_0 ;
  wire \read_data[13]_INST_0_i_13_n_0 ;
  wire \read_data[13]_INST_0_i_14_n_0 ;
  wire \read_data[13]_INST_0_i_15_n_0 ;
  wire \read_data[13]_INST_0_i_1_n_0 ;
  wire \read_data[13]_INST_0_i_2_n_0 ;
  wire \read_data[13]_INST_0_i_3_n_0 ;
  wire \read_data[13]_INST_0_i_4_n_0 ;
  wire \read_data[13]_INST_0_i_5_n_0 ;
  wire \read_data[13]_INST_0_i_6_n_0 ;
  wire \read_data[13]_INST_0_i_7_n_0 ;
  wire \read_data[13]_INST_0_i_8_n_0 ;
  wire \read_data[13]_INST_0_i_9_n_0 ;
  wire \read_data[14]_INST_0_i_10_n_0 ;
  wire \read_data[14]_INST_0_i_11_n_0 ;
  wire \read_data[14]_INST_0_i_12_n_0 ;
  wire \read_data[14]_INST_0_i_13_n_0 ;
  wire \read_data[14]_INST_0_i_1_n_0 ;
  wire \read_data[14]_INST_0_i_2_n_0 ;
  wire \read_data[14]_INST_0_i_3_n_0 ;
  wire \read_data[14]_INST_0_i_4_n_0 ;
  wire \read_data[14]_INST_0_i_5_n_0 ;
  wire \read_data[14]_INST_0_i_6_n_0 ;
  wire \read_data[14]_INST_0_i_7_n_0 ;
  wire \read_data[14]_INST_0_i_8_n_0 ;
  wire \read_data[14]_INST_0_i_9_n_0 ;
  wire \read_data[15]_INST_0_i_10_n_0 ;
  wire \read_data[15]_INST_0_i_11_n_0 ;
  wire \read_data[15]_INST_0_i_12_n_0 ;
  wire \read_data[15]_INST_0_i_13_n_0 ;
  wire \read_data[15]_INST_0_i_14_n_0 ;
  wire \read_data[15]_INST_0_i_15_n_0 ;
  wire \read_data[15]_INST_0_i_16_n_0 ;
  wire \read_data[15]_INST_0_i_1_n_0 ;
  wire \read_data[15]_INST_0_i_2_n_0 ;
  wire \read_data[15]_INST_0_i_3_n_0 ;
  wire \read_data[15]_INST_0_i_4_n_0 ;
  wire \read_data[15]_INST_0_i_5_n_0 ;
  wire \read_data[15]_INST_0_i_6_n_0 ;
  wire \read_data[15]_INST_0_i_7_n_0 ;
  wire \read_data[15]_INST_0_i_8_n_0 ;
  wire \read_data[15]_INST_0_i_9_n_0 ;
  wire \read_data[16]_INST_0_i_1_n_0 ;
  wire \read_data[16]_INST_0_i_2_n_0 ;
  wire \read_data[16]_INST_0_i_3_n_0 ;
  wire \read_data[16]_INST_0_i_4_n_0 ;
  wire \read_data[16]_INST_0_i_5_n_0 ;
  wire \read_data[16]_INST_0_i_6_n_0 ;
  wire \read_data[16]_INST_0_i_7_n_0 ;
  wire \read_data[16]_INST_0_i_8_n_0 ;
  wire \read_data[16]_INST_0_i_9_n_0 ;
  wire \read_data[17]_INST_0_i_10_n_0 ;
  wire \read_data[17]_INST_0_i_1_n_0 ;
  wire \read_data[17]_INST_0_i_2_n_0 ;
  wire \read_data[17]_INST_0_i_3_n_0 ;
  wire \read_data[17]_INST_0_i_4_n_0 ;
  wire \read_data[17]_INST_0_i_5_n_0 ;
  wire \read_data[17]_INST_0_i_6_n_0 ;
  wire \read_data[17]_INST_0_i_7_n_0 ;
  wire \read_data[17]_INST_0_i_8_n_0 ;
  wire \read_data[17]_INST_0_i_9_n_0 ;
  wire \read_data[18]_INST_0_i_1_n_0 ;
  wire \read_data[18]_INST_0_i_2_n_0 ;
  wire \read_data[18]_INST_0_i_3_n_0 ;
  wire \read_data[18]_INST_0_i_4_n_0 ;
  wire \read_data[18]_INST_0_i_5_n_0 ;
  wire \read_data[18]_INST_0_i_6_n_0 ;
  wire \read_data[18]_INST_0_i_7_n_0 ;
  wire \read_data[18]_INST_0_i_8_n_0 ;
  wire \read_data[19]_INST_0_i_1_n_0 ;
  wire \read_data[19]_INST_0_i_2_n_0 ;
  wire \read_data[19]_INST_0_i_3_n_0 ;
  wire \read_data[19]_INST_0_i_4_n_0 ;
  wire \read_data[19]_INST_0_i_5_n_0 ;
  wire \read_data[19]_INST_0_i_6_n_0 ;
  wire \read_data[19]_INST_0_i_7_n_0 ;
  wire \read_data[1]_INST_0_i_10_n_0 ;
  wire \read_data[1]_INST_0_i_1_n_0 ;
  wire \read_data[1]_INST_0_i_2_n_0 ;
  wire \read_data[1]_INST_0_i_3_n_0 ;
  wire \read_data[1]_INST_0_i_4_n_0 ;
  wire \read_data[1]_INST_0_i_5_n_0 ;
  wire \read_data[1]_INST_0_i_6_n_0 ;
  wire \read_data[1]_INST_0_i_7_n_0 ;
  wire \read_data[1]_INST_0_i_8_n_0 ;
  wire \read_data[1]_INST_0_i_9_n_0 ;
  wire \read_data[20]_INST_0_i_10_n_0 ;
  wire \read_data[20]_INST_0_i_1_n_0 ;
  wire \read_data[20]_INST_0_i_2_n_0 ;
  wire \read_data[20]_INST_0_i_3_n_0 ;
  wire \read_data[20]_INST_0_i_4_n_0 ;
  wire \read_data[20]_INST_0_i_5_n_0 ;
  wire \read_data[20]_INST_0_i_6_n_0 ;
  wire \read_data[20]_INST_0_i_7_n_0 ;
  wire \read_data[20]_INST_0_i_8_n_0 ;
  wire \read_data[20]_INST_0_i_9_n_0 ;
  wire \read_data[21]_INST_0_i_1_n_0 ;
  wire \read_data[21]_INST_0_i_2_n_0 ;
  wire \read_data[21]_INST_0_i_3_n_0 ;
  wire \read_data[21]_INST_0_i_4_n_0 ;
  wire \read_data[21]_INST_0_i_5_n_0 ;
  wire \read_data[21]_INST_0_i_6_n_0 ;
  wire \read_data[21]_INST_0_i_7_n_0 ;
  wire \read_data[21]_INST_0_i_8_n_0 ;
  wire \read_data[21]_INST_0_i_9_n_0 ;
  wire \read_data[22]_INST_0_i_1_n_0 ;
  wire \read_data[22]_INST_0_i_2_n_0 ;
  wire \read_data[22]_INST_0_i_3_n_0 ;
  wire \read_data[22]_INST_0_i_4_n_0 ;
  wire \read_data[22]_INST_0_i_5_n_0 ;
  wire \read_data[22]_INST_0_i_6_n_0 ;
  wire \read_data[22]_INST_0_i_7_n_0 ;
  wire \read_data[23]_INST_0_i_10_n_0 ;
  wire \read_data[23]_INST_0_i_11_n_0 ;
  wire \read_data[23]_INST_0_i_12_n_0 ;
  wire \read_data[23]_INST_0_i_1_n_0 ;
  wire \read_data[23]_INST_0_i_2_n_0 ;
  wire \read_data[23]_INST_0_i_3_n_0 ;
  wire \read_data[23]_INST_0_i_4_n_0 ;
  wire \read_data[23]_INST_0_i_5_n_0 ;
  wire \read_data[23]_INST_0_i_6_n_0 ;
  wire \read_data[23]_INST_0_i_7_n_0 ;
  wire \read_data[23]_INST_0_i_8_n_0 ;
  wire \read_data[23]_INST_0_i_9_n_0 ;
  wire \read_data[24]_INST_0_i_10_n_0 ;
  wire \read_data[24]_INST_0_i_11_n_0 ;
  wire \read_data[24]_INST_0_i_12_n_0 ;
  wire \read_data[24]_INST_0_i_13_n_0 ;
  wire \read_data[24]_INST_0_i_14_n_0 ;
  wire \read_data[24]_INST_0_i_15_n_0 ;
  wire \read_data[24]_INST_0_i_16_n_0 ;
  wire \read_data[24]_INST_0_i_1_n_0 ;
  wire \read_data[24]_INST_0_i_2_n_0 ;
  wire \read_data[24]_INST_0_i_3_n_0 ;
  wire \read_data[24]_INST_0_i_4_n_0 ;
  wire \read_data[24]_INST_0_i_5_n_0 ;
  wire \read_data[24]_INST_0_i_6_n_0 ;
  wire \read_data[24]_INST_0_i_7_n_0 ;
  wire \read_data[24]_INST_0_i_8_n_0 ;
  wire \read_data[24]_INST_0_i_9_n_0 ;
  wire \read_data[25]_INST_0_i_10_n_0 ;
  wire \read_data[25]_INST_0_i_11_n_0 ;
  wire \read_data[25]_INST_0_i_12_n_0 ;
  wire \read_data[25]_INST_0_i_13_n_0 ;
  wire \read_data[25]_INST_0_i_14_n_0 ;
  wire \read_data[25]_INST_0_i_15_n_0 ;
  wire \read_data[25]_INST_0_i_1_n_0 ;
  wire \read_data[25]_INST_0_i_2_n_0 ;
  wire \read_data[25]_INST_0_i_3_n_0 ;
  wire \read_data[25]_INST_0_i_4_n_0 ;
  wire \read_data[25]_INST_0_i_5_n_0 ;
  wire \read_data[25]_INST_0_i_6_n_0 ;
  wire \read_data[25]_INST_0_i_7_n_0 ;
  wire \read_data[25]_INST_0_i_8_n_0 ;
  wire \read_data[25]_INST_0_i_9_n_0 ;
  wire \read_data[26]_INST_0_i_1_n_0 ;
  wire \read_data[26]_INST_0_i_2_n_0 ;
  wire \read_data[26]_INST_0_i_3_n_0 ;
  wire \read_data[26]_INST_0_i_4_n_0 ;
  wire \read_data[26]_INST_0_i_5_n_0 ;
  wire \read_data[26]_INST_0_i_6_n_0 ;
  wire \read_data[26]_INST_0_i_7_n_0 ;
  wire \read_data[26]_INST_0_i_8_n_0 ;
  wire \read_data[27]_INST_0_i_10_n_0 ;
  wire \read_data[27]_INST_0_i_11_n_0 ;
  wire \read_data[27]_INST_0_i_12_n_0 ;
  wire \read_data[27]_INST_0_i_13_n_0 ;
  wire \read_data[27]_INST_0_i_1_n_0 ;
  wire \read_data[27]_INST_0_i_2_n_0 ;
  wire \read_data[27]_INST_0_i_3_n_0 ;
  wire \read_data[27]_INST_0_i_4_n_0 ;
  wire \read_data[27]_INST_0_i_5_n_0 ;
  wire \read_data[27]_INST_0_i_6_n_0 ;
  wire \read_data[27]_INST_0_i_7_n_0 ;
  wire \read_data[27]_INST_0_i_8_n_0 ;
  wire \read_data[27]_INST_0_i_9_n_0 ;
  wire \read_data[28]_INST_0_i_10_n_0 ;
  wire \read_data[28]_INST_0_i_11_n_0 ;
  wire \read_data[28]_INST_0_i_1_n_0 ;
  wire \read_data[28]_INST_0_i_2_n_0 ;
  wire \read_data[28]_INST_0_i_3_n_0 ;
  wire \read_data[28]_INST_0_i_4_n_0 ;
  wire \read_data[28]_INST_0_i_5_n_0 ;
  wire \read_data[28]_INST_0_i_6_n_0 ;
  wire \read_data[28]_INST_0_i_7_n_0 ;
  wire \read_data[28]_INST_0_i_8_n_0 ;
  wire \read_data[28]_INST_0_i_9_n_0 ;
  wire \read_data[29]_INST_0_i_10_n_0 ;
  wire \read_data[29]_INST_0_i_11_n_0 ;
  wire \read_data[29]_INST_0_i_12_n_0 ;
  wire \read_data[29]_INST_0_i_13_n_0 ;
  wire \read_data[29]_INST_0_i_14_n_0 ;
  wire \read_data[29]_INST_0_i_15_n_0 ;
  wire \read_data[29]_INST_0_i_1_n_0 ;
  wire \read_data[29]_INST_0_i_2_n_0 ;
  wire \read_data[29]_INST_0_i_3_n_0 ;
  wire \read_data[29]_INST_0_i_4_n_0 ;
  wire \read_data[29]_INST_0_i_5_n_0 ;
  wire \read_data[29]_INST_0_i_6_n_0 ;
  wire \read_data[29]_INST_0_i_7_n_0 ;
  wire \read_data[29]_INST_0_i_8_n_0 ;
  wire \read_data[29]_INST_0_i_9_n_0 ;
  wire \read_data[2]_INST_0_i_1_n_0 ;
  wire \read_data[2]_INST_0_i_2_n_0 ;
  wire \read_data[2]_INST_0_i_3_n_0 ;
  wire \read_data[2]_INST_0_i_4_n_0 ;
  wire \read_data[2]_INST_0_i_5_n_0 ;
  wire \read_data[2]_INST_0_i_6_n_0 ;
  wire \read_data[2]_INST_0_i_7_n_0 ;
  wire \read_data[30]_INST_0_i_10_n_0 ;
  wire \read_data[30]_INST_0_i_11_n_0 ;
  wire \read_data[30]_INST_0_i_12_n_0 ;
  wire \read_data[30]_INST_0_i_13_n_0 ;
  wire \read_data[30]_INST_0_i_1_n_0 ;
  wire \read_data[30]_INST_0_i_2_n_0 ;
  wire \read_data[30]_INST_0_i_3_n_0 ;
  wire \read_data[30]_INST_0_i_4_n_0 ;
  wire \read_data[30]_INST_0_i_5_n_0 ;
  wire \read_data[30]_INST_0_i_6_n_0 ;
  wire \read_data[30]_INST_0_i_7_n_0 ;
  wire \read_data[30]_INST_0_i_8_n_0 ;
  wire \read_data[30]_INST_0_i_9_n_0 ;
  wire \read_data[31]_INST_0_i_10_n_0 ;
  wire \read_data[31]_INST_0_i_11_n_0 ;
  wire \read_data[31]_INST_0_i_12_n_0 ;
  wire \read_data[31]_INST_0_i_13_n_0 ;
  wire \read_data[31]_INST_0_i_14_n_0 ;
  wire \read_data[31]_INST_0_i_15_n_0 ;
  wire \read_data[31]_INST_0_i_16_n_0 ;
  wire \read_data[31]_INST_0_i_1_n_0 ;
  wire \read_data[31]_INST_0_i_2_n_0 ;
  wire \read_data[31]_INST_0_i_3_n_0 ;
  wire \read_data[31]_INST_0_i_4_n_0 ;
  wire \read_data[31]_INST_0_i_5_n_0 ;
  wire \read_data[31]_INST_0_i_6_n_0 ;
  wire \read_data[31]_INST_0_i_7_n_0 ;
  wire \read_data[31]_INST_0_i_8_n_0 ;
  wire \read_data[31]_INST_0_i_9_n_0 ;
  wire \read_data[3]_INST_0_i_1_n_0 ;
  wire \read_data[3]_INST_0_i_2_n_0 ;
  wire \read_data[3]_INST_0_i_3_n_0 ;
  wire \read_data[3]_INST_0_i_4_n_0 ;
  wire \read_data[3]_INST_0_i_5_n_0 ;
  wire \read_data[3]_INST_0_i_6_n_0 ;
  wire \read_data[3]_INST_0_i_7_n_0 ;
  wire \read_data[4]_INST_0_i_1_n_0 ;
  wire \read_data[4]_INST_0_i_2_n_0 ;
  wire \read_data[4]_INST_0_i_3_n_0 ;
  wire \read_data[4]_INST_0_i_4_n_0 ;
  wire \read_data[4]_INST_0_i_5_n_0 ;
  wire \read_data[4]_INST_0_i_6_n_0 ;
  wire \read_data[4]_INST_0_i_7_n_0 ;
  wire \read_data[4]_INST_0_i_8_n_0 ;
  wire \read_data[4]_INST_0_i_9_n_0 ;
  wire \read_data[5]_INST_0_i_1_n_0 ;
  wire \read_data[5]_INST_0_i_2_n_0 ;
  wire \read_data[5]_INST_0_i_3_n_0 ;
  wire \read_data[5]_INST_0_i_4_n_0 ;
  wire \read_data[5]_INST_0_i_5_n_0 ;
  wire \read_data[5]_INST_0_i_6_n_0 ;
  wire \read_data[5]_INST_0_i_7_n_0 ;
  wire \read_data[5]_INST_0_i_8_n_0 ;
  wire \read_data[5]_INST_0_i_9_n_0 ;
  wire \read_data[6]_INST_0_i_1_n_0 ;
  wire \read_data[6]_INST_0_i_2_n_0 ;
  wire \read_data[6]_INST_0_i_3_n_0 ;
  wire \read_data[6]_INST_0_i_4_n_0 ;
  wire \read_data[6]_INST_0_i_5_n_0 ;
  wire \read_data[6]_INST_0_i_6_n_0 ;
  wire \read_data[6]_INST_0_i_7_n_0 ;
  wire \read_data[7]_INST_0_i_1_n_0 ;
  wire \read_data[7]_INST_0_i_2_n_0 ;
  wire \read_data[7]_INST_0_i_3_n_0 ;
  wire \read_data[7]_INST_0_i_4_n_0 ;
  wire \read_data[7]_INST_0_i_5_n_0 ;
  wire \read_data[7]_INST_0_i_6_n_0 ;
  wire \read_data[7]_INST_0_i_7_n_0 ;
  wire \read_data[8]_INST_0_i_10_n_0 ;
  wire \read_data[8]_INST_0_i_11_n_0 ;
  wire \read_data[8]_INST_0_i_12_n_0 ;
  wire \read_data[8]_INST_0_i_13_n_0 ;
  wire \read_data[8]_INST_0_i_14_n_0 ;
  wire \read_data[8]_INST_0_i_15_n_0 ;
  wire \read_data[8]_INST_0_i_16_n_0 ;
  wire \read_data[8]_INST_0_i_1_n_0 ;
  wire \read_data[8]_INST_0_i_2_n_0 ;
  wire \read_data[8]_INST_0_i_3_n_0 ;
  wire \read_data[8]_INST_0_i_4_n_0 ;
  wire \read_data[8]_INST_0_i_5_n_0 ;
  wire \read_data[8]_INST_0_i_6_n_0 ;
  wire \read_data[8]_INST_0_i_7_n_0 ;
  wire \read_data[8]_INST_0_i_8_n_0 ;
  wire \read_data[8]_INST_0_i_9_n_0 ;
  wire \read_data[9]_INST_0_i_10_n_0 ;
  wire \read_data[9]_INST_0_i_11_n_0 ;
  wire \read_data[9]_INST_0_i_12_n_0 ;
  wire \read_data[9]_INST_0_i_13_n_0 ;
  wire \read_data[9]_INST_0_i_14_n_0 ;
  wire \read_data[9]_INST_0_i_15_n_0 ;
  wire \read_data[9]_INST_0_i_1_n_0 ;
  wire \read_data[9]_INST_0_i_2_n_0 ;
  wire \read_data[9]_INST_0_i_3_n_0 ;
  wire \read_data[9]_INST_0_i_4_n_0 ;
  wire \read_data[9]_INST_0_i_5_n_0 ;
  wire \read_data[9]_INST_0_i_6_n_0 ;
  wire \read_data[9]_INST_0_i_7_n_0 ;
  wire \read_data[9]_INST_0_i_8_n_0 ;
  wire \read_data[9]_INST_0_i_9_n_0 ;

  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[0]_INST_0 
       (.I0(\read_data[0]_INST_0_i_1_n_0 ),
        .I1(addr[8]),
        .I2(\read_data[0]_INST_0_i_2_n_0 ),
        .I3(addr[7]),
        .I4(\read_data[0]_INST_0_i_3_n_0 ),
        .O(read_data[0]));
  MUXF7 \read_data[0]_INST_0_i_1 
       (.I0(\read_data[0]_INST_0_i_4_n_0 ),
        .I1(\read_data[0]_INST_0_i_5_n_0 ),
        .O(\read_data[0]_INST_0_i_1_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[0]_INST_0_i_2 
       (.I0(\read_data[0]_INST_0_i_6_n_0 ),
        .I1(\read_data[0]_INST_0_i_7_n_0 ),
        .O(\read_data[0]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[0]_INST_0_i_3 
       (.I0(\read_data[0]_INST_0_i_8_n_0 ),
        .I1(\read_data[0]_INST_0_i_9_n_0 ),
        .O(\read_data[0]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h0000FFFF80FF0000)) 
    \read_data[0]_INST_0_i_4 
       (.I0(addr[3]),
        .I1(addr[4]),
        .I2(addr[6]),
        .I3(addr[5]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0777000074440000)) 
    \read_data[0]_INST_0_i_5 
       (.I0(addr[6]),
        .I1(addr[0]),
        .I2(addr[3]),
        .I3(addr[4]),
        .I4(addr[2]),
        .I5(addr[5]),
        .O(\read_data[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4002212022220000)) 
    \read_data[0]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[4]),
        .O(\read_data[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h83080E000E750E00)) 
    \read_data[0]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(addr[5]),
        .I2(addr[2]),
        .I3(addr[6]),
        .I4(addr[4]),
        .I5(addr[3]),
        .O(\read_data[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00010800155515D5)) 
    \read_data[0]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[4]),
        .I3(addr[5]),
        .I4(addr[3]),
        .I5(addr[2]),
        .O(\read_data[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000401041)) 
    \read_data[0]_INST_0_i_9 
       (.I0(addr[6]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[0]),
        .O(\read_data[0]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[10]_INST_0 
       (.I0(\read_data[10]_INST_0_i_1_n_0 ),
        .I1(\read_data[15]_INST_0_i_2_n_0 ),
        .I2(\read_data[10]_INST_0_i_2_n_0 ),
        .I3(\read_data[15]_INST_0_i_4_n_0 ),
        .I4(\read_data[10]_INST_0_i_3_n_0 ),
        .O(read_data[10]));
  LUT6 #(
    .INIT(64'h0CFF05F00CF005F0)) 
    \read_data[10]_INST_0_i_1 
       (.I0(addr[2]),
        .I1(\read_data[12]_INST_0_i_4_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[13]_INST_0_i_8_n_0 ),
        .O(\read_data[10]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[10]_INST_0_i_2 
       (.I0(\read_data[10]_INST_0_i_4_n_0 ),
        .I1(\read_data[11]_INST_0_i_7_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[12]_INST_0_i_7_n_0 ),
        .I5(\read_data[10]_INST_0_i_5_n_0 ),
        .O(\read_data[10]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hCB0BC808)) 
    \read_data[10]_INST_0_i_3 
       (.I0(\read_data[10]_INST_0_i_6_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[10]_INST_0_i_7_n_0 ),
        .I4(\read_data[10]_INST_0_i_8_n_0 ),
        .O(\read_data[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEBC3C3C3D7FFBFFD)) 
    \read_data[10]_INST_0_i_4 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[10]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02800000557FEA82)) 
    \read_data[10]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[10]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFEA00004142416B)) 
    \read_data[10]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[10]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000056AA5557AAA8)) 
    \read_data[10]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[10]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0014028028001400)) 
    \read_data[10]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[11]_INST_0 
       (.I0(\read_data[11]_INST_0_i_1_n_0 ),
        .I1(\read_data[11]_INST_0_i_2_n_0 ),
        .I2(\read_data[15]_INST_0_i_2_n_0 ),
        .I3(\read_data[11]_INST_0_i_3_n_0 ),
        .I4(\read_data[15]_INST_0_i_4_n_0 ),
        .I5(\read_data[11]_INST_0_i_4_n_0 ),
        .O(read_data[11]));
  LUT5 #(
    .INIT(32'hFCAF0CA0)) 
    \read_data[11]_INST_0_i_1 
       (.I0(\read_data[13]_INST_0_i_5_n_0 ),
        .I1(\read_data[11]_INST_0_i_5_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[11]_INST_0_i_6_n_0 ),
        .O(\read_data[11]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000006A6A000000)) 
    \read_data[11]_INST_0_i_10 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[11]_INST_0_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'h01101010)) 
    \read_data[11]_INST_0_i_11 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[2]),
        .I3(addr[0]),
        .I4(addr[1]),
        .O(\read_data[11]_INST_0_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \read_data[11]_INST_0_i_12 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .O(\read_data[11]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h9000000300030003)) 
    \read_data[11]_INST_0_i_13 
       (.I0(addr[4]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[0]),
        .I5(addr[1]),
        .O(\read_data[11]_INST_0_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \read_data[11]_INST_0_i_2 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .O(\read_data[11]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFCAF0CA0)) 
    \read_data[11]_INST_0_i_3 
       (.I0(\read_data[13]_INST_0_i_5_n_0 ),
        .I1(\read_data[11]_INST_0_i_7_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[11]_INST_0_i_6_n_0 ),
        .O(\read_data[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hC303C000C808C808)) 
    \read_data[11]_INST_0_i_4 
       (.I0(\read_data[11]_INST_0_i_8_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[11]_INST_0_i_9_n_0 ),
        .I4(\read_data[11]_INST_0_i_10_n_0 ),
        .I5(\read_data[15]_INST_0_i_9_n_0 ),
        .O(\read_data[11]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD7FFFFFFFFFFEBC3)) 
    \read_data[11]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[11]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB08000000000B080)) 
    \read_data[11]_INST_0_i_6 
       (.I0(\read_data[11]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[11]_INST_0_i_12_n_0 ),
        .I3(\read_data[11]_INST_0_i_13_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[15]_INST_0_i_6_n_0 ),
        .O(\read_data[11]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h16BC3C3C7D7FEA82)) 
    \read_data[11]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[11]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0015EA0000000000)) 
    \read_data[11]_INST_0_i_8 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0155A8005557AAA8)) 
    \read_data[11]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[11]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[12]_INST_0 
       (.I0(\read_data[12]_INST_0_i_1_n_0 ),
        .I1(\read_data[15]_INST_0_i_2_n_0 ),
        .I2(\read_data[12]_INST_0_i_2_n_0 ),
        .I3(\read_data[15]_INST_0_i_4_n_0 ),
        .I4(\read_data[12]_INST_0_i_3_n_0 ),
        .O(read_data[12]));
  LUT6 #(
    .INIT(64'h0C0F05000C000500)) 
    \read_data[12]_INST_0_i_1 
       (.I0(addr[2]),
        .I1(\read_data[12]_INST_0_i_4_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[13]_INST_0_i_8_n_0 ),
        .O(\read_data[12]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000001AAA80000)) 
    \read_data[12]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0015800028001400)) 
    \read_data[12]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[12]_INST_0_i_2 
       (.I0(\read_data[12]_INST_0_i_5_n_0 ),
        .I1(\read_data[12]_INST_0_i_6_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[12]_INST_0_i_7_n_0 ),
        .I5(\read_data[13]_INST_0_i_14_n_0 ),
        .O(\read_data[12]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[12]_INST_0_i_3 
       (.I0(\read_data[12]_INST_0_i_8_n_0 ),
        .I1(\read_data[12]_INST_0_i_9_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[12]_INST_0_i_10_n_0 ),
        .I5(\read_data[12]_INST_0_i_11_n_0 ),
        .O(\read_data[12]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEBBBC333C333C333)) 
    \read_data[12]_INST_0_i_4 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h143C3C3C28000000)) 
    \read_data[12]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h96BC3C3C7D7FFFD7)) 
    \read_data[12]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4143C3C382800000)) 
    \read_data[12]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0004040444545440)) 
    \read_data[12]_INST_0_i_8 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[15]_INST_0_i_16_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFEBFFFFFAAA9BEBD)) 
    \read_data[12]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[12]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[13]_INST_0 
       (.I0(\read_data[13]_INST_0_i_1_n_0 ),
        .I1(\read_data[13]_INST_0_i_2_n_0 ),
        .I2(\read_data[15]_INST_0_i_2_n_0 ),
        .I3(\read_data[13]_INST_0_i_3_n_0 ),
        .I4(\read_data[15]_INST_0_i_4_n_0 ),
        .I5(\read_data[13]_INST_0_i_4_n_0 ),
        .O(read_data[13]));
  LUT5 #(
    .INIT(32'hFB3BF838)) 
    \read_data[13]_INST_0_i_1 
       (.I0(\read_data[13]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[13]_INST_0_i_6_n_0 ),
        .I4(\read_data[13]_INST_0_i_7_n_0 ),
        .O(\read_data[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h294003C016BC6802)) 
    \read_data[13]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[13]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000444444440)) 
    \read_data[13]_INST_0_i_11 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[15]_INST_0_i_16_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[13]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7EAA000055564142)) 
    \read_data[13]_INST_0_i_12 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8014001580019401)) 
    \read_data[13]_INST_0_i_13 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[13]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000110000000)) 
    \read_data[13]_INST_0_i_14 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[15]_INST_0_i_16_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[13]_INST_0_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \read_data[13]_INST_0_i_15 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .O(\read_data[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD555C444C444C444)) 
    \read_data[13]_INST_0_i_2 
       (.I0(addr[0]),
        .I1(addr[1]),
        .I2(\read_data[13]_INST_0_i_8_n_0 ),
        .I3(\read_data[15]_INST_0_i_9_n_0 ),
        .I4(addr[3]),
        .I5(addr[2]),
        .O(\read_data[13]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3B3BFB3B3838F838)) 
    \read_data[13]_INST_0_i_3 
       (.I0(\read_data[13]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[13]_INST_0_i_9_n_0 ),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[13]_INST_0_i_10_n_0 ),
        .O(\read_data[13]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[13]_INST_0_i_4 
       (.I0(\read_data[13]_INST_0_i_11_n_0 ),
        .I1(\read_data[13]_INST_0_i_12_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[13]_INST_0_i_13_n_0 ),
        .I5(\read_data[13]_INST_0_i_14_n_0 ),
        .O(\read_data[13]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h11155444)) 
    \read_data[13]_INST_0_i_5 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[13]_INST_0_i_15_n_0 ),
        .I4(addr[4]),
        .O(\read_data[13]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2A80000041438280)) 
    \read_data[13]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[13]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h3D403FC03EBC3C00)) 
    \read_data[13]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[13]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0880808080808080)) 
    \read_data[13]_INST_0_i_8 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0015959595800000)) 
    \read_data[13]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[13]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[14]_INST_0 
       (.I0(\read_data[14]_INST_0_i_1_n_0 ),
        .I1(\read_data[14]_INST_0_i_2_n_0 ),
        .I2(\read_data[15]_INST_0_i_2_n_0 ),
        .I3(\read_data[14]_INST_0_i_3_n_0 ),
        .I4(\read_data[15]_INST_0_i_4_n_0 ),
        .I5(\read_data[14]_INST_0_i_4_n_0 ),
        .O(read_data[14]));
  LUT5 #(
    .INIT(32'hEB2BE828)) 
    \read_data[14]_INST_0_i_1 
       (.I0(\read_data[14]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[14]_INST_0_i_6_n_0 ),
        .I4(\read_data[14]_INST_0_i_7_n_0 ),
        .O(\read_data[14]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8015FFEA15959595)) 
    \read_data[14]_INST_0_i_10 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[14]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0014014180001400)) 
    \read_data[14]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[14]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0080808080000000)) 
    \read_data[14]_INST_0_i_12 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h6A7FFFFFFF958000)) 
    \read_data[14]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[14]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFF00000000009090)) 
    \read_data[14]_INST_0_i_2 
       (.I0(addr[4]),
        .I1(addr[3]),
        .I2(addr[2]),
        .I3(\read_data[14]_INST_0_i_8_n_0 ),
        .I4(addr[1]),
        .I5(addr[0]),
        .O(\read_data[14]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h2B2BEB2B2828E828)) 
    \read_data[14]_INST_0_i_3 
       (.I0(\read_data[14]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[14]_INST_0_i_9_n_0 ),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[14]_INST_0_i_7_n_0 ),
        .O(\read_data[14]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF0000044)) 
    \read_data[14]_INST_0_i_4 
       (.I0(\read_data[15]_INST_0_i_9_n_0 ),
        .I1(\read_data[14]_INST_0_i_10_n_0 ),
        .I2(\read_data[14]_INST_0_i_11_n_0 ),
        .I3(addr[1]),
        .I4(addr[0]),
        .O(\read_data[14]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBF0F0BB88F0F088)) 
    \read_data[14]_INST_0_i_5 
       (.I0(\read_data[14]_INST_0_i_12_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[8]_INST_0_i_5_n_0 ),
        .I3(\read_data[15]_INST_0_i_6_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[14]_INST_0_i_13_n_0 ),
        .O(\read_data[14]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hC003C003D403E803)) 
    \read_data[14]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[14]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2801828197C06AAA)) 
    \read_data[14]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[14]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEA83C003C003C003)) 
    \read_data[14]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0015EA15EA158000)) 
    \read_data[14]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[14]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[15]_INST_0 
       (.I0(\read_data[15]_INST_0_i_1_n_0 ),
        .I1(\read_data[15]_INST_0_i_2_n_0 ),
        .I2(\read_data[15]_INST_0_i_3_n_0 ),
        .I3(\read_data[15]_INST_0_i_4_n_0 ),
        .I4(\read_data[15]_INST_0_i_5_n_0 ),
        .O(read_data[15]));
  LUT6 #(
    .INIT(64'h8414149494040484)) 
    \read_data[15]_INST_0_i_1 
       (.I0(addr[0]),
        .I1(addr[1]),
        .I2(addr[2]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[15]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4143828015558000)) 
    \read_data[15]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[15]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0015FFEA00001580)) 
    \read_data[15]_INST_0_i_11 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[15]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0012121212000000)) 
    \read_data[15]_INST_0_i_12 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h1580000000006A00)) 
    \read_data[15]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[15]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hC1114333C333C333)) 
    \read_data[15]_INST_0_i_14 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h1804040404848484)) 
    \read_data[15]_INST_0_i_15 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[15]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \read_data[15]_INST_0_i_16 
       (.I0(addr[1]),
        .I1(addr[0]),
        .O(\read_data[15]_INST_0_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \read_data[15]_INST_0_i_2 
       (.I0(addr[6]),
        .I1(\read_data[15]_INST_0_i_6_n_0 ),
        .I2(addr[7]),
        .I3(addr[8]),
        .O(\read_data[15]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h2B2BEB2B2828E828)) 
    \read_data[15]_INST_0_i_3 
       (.I0(\read_data[15]_INST_0_i_7_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[15]_INST_0_i_8_n_0 ),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[15]_INST_0_i_10_n_0 ),
        .O(\read_data[15]_INST_0_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \read_data[15]_INST_0_i_4 
       (.I0(\read_data[15]_INST_0_i_6_n_0 ),
        .I1(addr[6]),
        .I2(addr[7]),
        .O(\read_data[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hC000C0000B0B0808)) 
    \read_data[15]_INST_0_i_5 
       (.I0(\read_data[15]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[15]_INST_0_i_12_n_0 ),
        .I4(\read_data[15]_INST_0_i_13_n_0 ),
        .I5(\read_data[15]_INST_0_i_9_n_0 ),
        .O(\read_data[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \read_data[15]_INST_0_i_6 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC0C0AFA0AFA0C0C0)) 
    \read_data[15]_INST_0_i_7 
       (.I0(\read_data[15]_INST_0_i_14_n_0 ),
        .I1(\read_data[15]_INST_0_i_15_n_0 ),
        .I2(addr[0]),
        .I3(\read_data[9]_INST_0_i_8_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[15]_INST_0_i_6_n_0 ),
        .O(\read_data[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0015FFEA00158000)) 
    \read_data[15]_INST_0_i_8 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[15]_INST_0_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \read_data[15]_INST_0_i_9 
       (.I0(\read_data[15]_INST_0_i_6_n_0 ),
        .I1(addr[6]),
        .O(\read_data[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[16]_INST_0 
       (.I0(\read_data[16]_INST_0_i_1_n_0 ),
        .I1(\read_data[23]_INST_0_i_1_n_0 ),
        .I2(\read_data[16]_INST_0_i_2_n_0 ),
        .I3(\read_data[18]_INST_0_i_3_n_0 ),
        .I4(\read_data[16]_INST_0_i_3_n_0 ),
        .O(read_data[16]));
  MUXF7 \read_data[16]_INST_0_i_1 
       (.I0(\read_data[16]_INST_0_i_4_n_0 ),
        .I1(\read_data[16]_INST_0_i_5_n_0 ),
        .O(\read_data[16]_INST_0_i_1_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[16]_INST_0_i_2 
       (.I0(\read_data[16]_INST_0_i_6_n_0 ),
        .I1(\read_data[16]_INST_0_i_7_n_0 ),
        .O(\read_data[16]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[16]_INST_0_i_3 
       (.I0(\read_data[16]_INST_0_i_8_n_0 ),
        .I1(\read_data[16]_INST_0_i_9_n_0 ),
        .O(\read_data[16]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h0777000074440000)) 
    \read_data[16]_INST_0_i_4 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[23]_INST_0_i_12_n_0 ),
        .O(\read_data[16]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFF80FF0000)) 
    \read_data[16]_INST_0_i_5 
       (.I0(\read_data[23]_INST_0_i_10_n_0 ),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[20]_INST_0_i_7_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(addr[0]),
        .I5(\read_data[23]_INST_0_i_11_n_0 ),
        .O(\read_data[16]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h83080E000E750E00)) 
    \read_data[16]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_12_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[20]_INST_0_i_7_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[23]_INST_0_i_10_n_0 ),
        .O(\read_data[16]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4002212022220000)) 
    \read_data[16]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[16]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000401041)) 
    \read_data[16]_INST_0_i_8 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(addr[0]),
        .O(\read_data[16]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00010800155515D5)) 
    \read_data[16]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[23]_INST_0_i_11_n_0 ),
        .O(\read_data[16]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[17]_INST_0 
       (.I0(\read_data[17]_INST_0_i_1_n_0 ),
        .I1(\read_data[23]_INST_0_i_1_n_0 ),
        .I2(\read_data[17]_INST_0_i_2_n_0 ),
        .I3(\read_data[18]_INST_0_i_3_n_0 ),
        .I4(\read_data[17]_INST_0_i_3_n_0 ),
        .O(read_data[17]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \read_data[17]_INST_0_i_1 
       (.I0(\read_data[17]_INST_0_i_4_n_0 ),
        .I1(\read_data[18]_INST_0_i_3_n_0 ),
        .I2(\read_data[17]_INST_0_i_5_n_0 ),
        .I3(addr[1]),
        .I4(\read_data[17]_INST_0_i_6_n_0 ),
        .O(\read_data[17]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h110C31C704114406)) 
    \read_data[17]_INST_0_i_10 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[23]_INST_0_i_11_n_0 ),
        .O(\read_data[17]_INST_0_i_10_n_0 ));
  MUXF7 \read_data[17]_INST_0_i_2 
       (.I0(\read_data[17]_INST_0_i_7_n_0 ),
        .I1(\read_data[17]_INST_0_i_8_n_0 ),
        .O(\read_data[17]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[17]_INST_0_i_3 
       (.I0(\read_data[17]_INST_0_i_9_n_0 ),
        .I1(\read_data[17]_INST_0_i_10_n_0 ),
        .O(\read_data[17]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'hFCCC0000CFFF0400)) 
    \read_data[17]_INST_0_i_4 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[23]_INST_0_i_12_n_0 ),
        .O(\read_data[17]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5111111100000000)) 
    \read_data[17]_INST_0_i_5 
       (.I0(\read_data[23]_INST_0_i_11_n_0 ),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(addr[0]),
        .O(\read_data[17]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3C282828283C3C3C)) 
    \read_data[17]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[17]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC002388E000088CC)) 
    \read_data[17]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[17]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h2A00AA0080008408)) 
    \read_data[17]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[17]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000401)) 
    \read_data[17]_INST_0_i_9 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(addr[0]),
        .O(\read_data[17]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[18]_INST_0 
       (.I0(\read_data[18]_INST_0_i_1_n_0 ),
        .I1(\read_data[23]_INST_0_i_1_n_0 ),
        .I2(\read_data[18]_INST_0_i_2_n_0 ),
        .I3(\read_data[18]_INST_0_i_3_n_0 ),
        .I4(\read_data[18]_INST_0_i_4_n_0 ),
        .O(read_data[18]));
  LUT6 #(
    .INIT(64'h80FF800000FF00FF)) 
    \read_data[18]_INST_0_i_1 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(\read_data[20]_INST_0_i_8_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(addr[1]),
        .I4(\read_data[20]_INST_0_i_10_n_0 ),
        .I5(addr[0]),
        .O(\read_data[18]_INST_0_i_1_n_0 ));
  MUXF7 \read_data[18]_INST_0_i_2 
       (.I0(\read_data[18]_INST_0_i_5_n_0 ),
        .I1(\read_data[18]_INST_0_i_6_n_0 ),
        .O(\read_data[18]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \read_data[18]_INST_0_i_3 
       (.I0(\read_data[23]_INST_0_i_4_n_0 ),
        .I1(addr[7]),
        .O(\read_data[18]_INST_0_i_3_n_0 ));
  MUXF7 \read_data[18]_INST_0_i_4 
       (.I0(\read_data[18]_INST_0_i_7_n_0 ),
        .I1(\read_data[18]_INST_0_i_8_n_0 ),
        .O(\read_data[18]_INST_0_i_4_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h6DB7B796B795B795)) 
    \read_data[18]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[18]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0220966622006644)) 
    \read_data[18]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[18]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAA00731)) 
    \read_data[18]_INST_0_i_7 
       (.I0(\read_data[23]_INST_0_i_12_n_0 ),
        .I1(\read_data[23]_INST_0_i_11_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[20]_INST_0_i_7_n_0 ),
        .I5(addr[0]),
        .O(\read_data[18]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h2001191115D46000)) 
    \read_data[18]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[23]_INST_0_i_12_n_0 ),
        .O(\read_data[18]_INST_0_i_8_n_0 ));
  MUXF7 \read_data[19]_INST_0 
       (.I0(\read_data[19]_INST_0_i_1_n_0 ),
        .I1(\read_data[19]_INST_0_i_2_n_0 ),
        .O(read_data[19]),
        .S(\read_data[23]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[19]_INST_0_i_1 
       (.I0(\read_data[19]_INST_0_i_3_n_0 ),
        .I1(\read_data[19]_INST_0_i_4_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(\read_data[19]_INST_0_i_5_n_0 ),
        .I4(addr[1]),
        .I5(\read_data[19]_INST_0_i_6_n_0 ),
        .O(\read_data[19]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA0A0A0A0C0CFC0C0)) 
    \read_data[19]_INST_0_i_2 
       (.I0(\read_data[19]_INST_0_i_3_n_0 ),
        .I1(\read_data[19]_INST_0_i_7_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(addr[2]),
        .I4(addr[0]),
        .I5(addr[1]),
        .O(\read_data[19]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000408)) 
    \read_data[19]_INST_0_i_3 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[19]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h488888888FF0F7F0)) 
    \read_data[19]_INST_0_i_4 
       (.I0(\read_data[23]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[19]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00011D55D1100000)) 
    \read_data[19]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[23]_INST_0_i_12_n_0 ),
        .O(\read_data[19]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000040)) 
    \read_data[19]_INST_0_i_6 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(addr[0]),
        .O(\read_data[19]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4CCCCCCCCFF4F7F4)) 
    \read_data[19]_INST_0_i_7 
       (.I0(\read_data[23]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[19]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[1]_INST_0 
       (.I0(\read_data[1]_INST_0_i_1_n_0 ),
        .I1(addr[8]),
        .I2(\read_data[1]_INST_0_i_2_n_0 ),
        .I3(addr[7]),
        .I4(\read_data[1]_INST_0_i_3_n_0 ),
        .O(read_data[1]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \read_data[1]_INST_0_i_1 
       (.I0(\read_data[1]_INST_0_i_4_n_0 ),
        .I1(addr[7]),
        .I2(\read_data[1]_INST_0_i_5_n_0 ),
        .I3(addr[1]),
        .I4(\read_data[1]_INST_0_i_6_n_0 ),
        .O(\read_data[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000401)) 
    \read_data[1]_INST_0_i_10 
       (.I0(addr[6]),
        .I1(addr[4]),
        .I2(addr[5]),
        .I3(addr[2]),
        .I4(addr[3]),
        .I5(addr[0]),
        .O(\read_data[1]_INST_0_i_10_n_0 ));
  MUXF7 \read_data[1]_INST_0_i_2 
       (.I0(\read_data[1]_INST_0_i_7_n_0 ),
        .I1(\read_data[1]_INST_0_i_8_n_0 ),
        .O(\read_data[1]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[1]_INST_0_i_3 
       (.I0(\read_data[1]_INST_0_i_9_n_0 ),
        .I1(\read_data[1]_INST_0_i_10_n_0 ),
        .O(\read_data[1]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'hFCCC0000CFFF0400)) 
    \read_data[1]_INST_0_i_4 
       (.I0(addr[6]),
        .I1(addr[0]),
        .I2(addr[3]),
        .I3(addr[4]),
        .I4(addr[2]),
        .I5(addr[5]),
        .O(\read_data[1]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEA00BF00)) 
    \read_data[1]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(addr[3]),
        .I2(addr[4]),
        .I3(addr[2]),
        .I4(addr[5]),
        .O(\read_data[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5111111100000000)) 
    \read_data[1]_INST_0_i_6 
       (.I0(addr[2]),
        .I1(addr[6]),
        .I2(addr[4]),
        .I3(addr[5]),
        .I4(addr[3]),
        .I5(addr[0]),
        .O(\read_data[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2A00AA0080008408)) 
    \read_data[1]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(addr[4]),
        .I2(addr[5]),
        .I3(addr[2]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hC002388E000088CC)) 
    \read_data[1]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[5]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h110C31C704114406)) 
    \read_data[1]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[4]),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[2]),
        .O(\read_data[1]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[20]_INST_0 
       (.I0(\read_data[20]_INST_0_i_1_n_0 ),
        .I1(\read_data[20]_INST_0_i_2_n_0 ),
        .O(read_data[20]),
        .S(\read_data[23]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[20]_INST_0_i_1 
       (.I0(\read_data[20]_INST_0_i_3_n_0 ),
        .I1(\read_data[20]_INST_0_i_4_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(\read_data[20]_INST_0_i_5_n_0 ),
        .I4(addr[1]),
        .I5(\read_data[20]_INST_0_i_6_n_0 ),
        .O(\read_data[20]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEBC3C3C3C3C3C3C3)) 
    \read_data[20]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[20]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h80FF800000000000)) 
    \read_data[20]_INST_0_i_2 
       (.I0(\read_data[20]_INST_0_i_7_n_0 ),
        .I1(\read_data[20]_INST_0_i_8_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(addr[1]),
        .I4(\read_data[20]_INST_0_i_10_n_0 ),
        .I5(addr[0]),
        .O(\read_data[20]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000144600004444)) 
    \read_data[20]_INST_0_i_3 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[20]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h3E82EC22EE22EE22)) 
    \read_data[20]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[20]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3010100002008084)) 
    \read_data[20]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[20]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA2AAAAE4746A)) 
    \read_data[20]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_12_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[20]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \read_data[20]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[20]_INST_0_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'h2888)) 
    \read_data[20]_INST_0_i_8 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[2]),
        .I3(addr[1]),
        .O(\read_data[20]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h7F80)) 
    \read_data[20]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[3]),
        .I3(addr[4]),
        .O(\read_data[20]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[21]_INST_0 
       (.I0(\read_data[21]_INST_0_i_1_n_0 ),
        .I1(\read_data[21]_INST_0_i_2_n_0 ),
        .O(read_data[21]),
        .S(\read_data[23]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8FFFFBBB80000)) 
    \read_data[21]_INST_0_i_1 
       (.I0(\read_data[21]_INST_0_i_3_n_0 ),
        .I1(addr[1]),
        .I2(\read_data[21]_INST_0_i_4_n_0 ),
        .I3(addr[0]),
        .I4(\read_data[18]_INST_0_i_3_n_0 ),
        .I5(\read_data[21]_INST_0_i_5_n_0 ),
        .O(\read_data[21]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0FFFFAFA0C0C0)) 
    \read_data[21]_INST_0_i_2 
       (.I0(\read_data[21]_INST_0_i_6_n_0 ),
        .I1(\read_data[21]_INST_0_i_4_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(\read_data[21]_INST_0_i_7_n_0 ),
        .I4(addr[1]),
        .I5(addr[0]),
        .O(\read_data[21]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8222000029909290)) 
    \read_data[21]_INST_0_i_3 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_11_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[21]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1115151554444444)) 
    \read_data[21]_INST_0_i_4 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[21]_INST_0_i_4_n_0 ));
  MUXF7 \read_data[21]_INST_0_i_5 
       (.I0(\read_data[21]_INST_0_i_8_n_0 ),
        .I1(\read_data[21]_INST_0_i_9_n_0 ),
        .O(\read_data[21]_INST_0_i_5_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'hE2A2A0A061919080)) 
    \read_data[21]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[20]_INST_0_i_9_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[23]_INST_0_i_11_n_0 ),
        .O(\read_data[21]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB888000088880000)) 
    \read_data[21]_INST_0_i_7 
       (.I0(\read_data[23]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[21]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88888000000ECEC0)) 
    \read_data[21]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_12_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[21]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200411045)) 
    \read_data[21]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[21]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[22]_INST_0 
       (.I0(\read_data[22]_INST_0_i_1_n_0 ),
        .I1(\read_data[22]_INST_0_i_2_n_0 ),
        .O(read_data[22]),
        .S(\read_data[23]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFA0C0C0)) 
    \read_data[22]_INST_0_i_1 
       (.I0(\read_data[22]_INST_0_i_3_n_0 ),
        .I1(\read_data[22]_INST_0_i_4_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(\read_data[22]_INST_0_i_5_n_0 ),
        .I4(addr[1]),
        .O(\read_data[22]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFA0C0C0)) 
    \read_data[22]_INST_0_i_2 
       (.I0(\read_data[22]_INST_0_i_6_n_0 ),
        .I1(\read_data[22]_INST_0_i_4_n_0 ),
        .I2(\read_data[18]_INST_0_i_3_n_0 ),
        .I3(\read_data[22]_INST_0_i_7_n_0 ),
        .I4(addr[1]),
        .O(\read_data[22]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h820000222E1BE010)) 
    \read_data[22]_INST_0_i_3 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_11_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[22]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h3E02EC22EE22CC00)) 
    \read_data[22]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[22]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0002002226201066)) 
    \read_data[22]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[22]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8330002022A05D7D)) 
    \read_data[22]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[23]_INST_0_i_12_n_0 ),
        .I4(\read_data[23]_INST_0_i_10_n_0 ),
        .I5(\read_data[23]_INST_0_i_11_n_0 ),
        .O(\read_data[22]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE0A040000A0A5555)) 
    \read_data[22]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_12_n_0 ),
        .I2(\read_data[20]_INST_0_i_9_n_0 ),
        .I3(\read_data[20]_INST_0_i_7_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[23]_INST_0_i_10_n_0 ),
        .O(\read_data[22]_INST_0_i_7_n_0 ));
  MUXF7 \read_data[23]_INST_0 
       (.I0(\read_data[23]_INST_0_i_2_n_0 ),
        .I1(\read_data[23]_INST_0_i_3_n_0 ),
        .O(read_data[23]),
        .S(\read_data[23]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \read_data[23]_INST_0_i_1 
       (.I0(\read_data[23]_INST_0_i_4_n_0 ),
        .I1(addr[7]),
        .I2(addr[8]),
        .O(\read_data[23]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \read_data[23]_INST_0_i_10 
       (.I0(addr[1]),
        .I1(addr[2]),
        .I2(addr[3]),
        .O(\read_data[23]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \read_data[23]_INST_0_i_11 
       (.I0(addr[1]),
        .I1(addr[2]),
        .O(\read_data[23]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \read_data[23]_INST_0_i_12 
       (.I0(addr[3]),
        .I1(addr[1]),
        .I2(addr[2]),
        .I3(addr[4]),
        .I4(addr[5]),
        .O(\read_data[23]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888B8BBB888)) 
    \read_data[23]_INST_0_i_2 
       (.I0(\read_data[23]_INST_0_i_5_n_0 ),
        .I1(\read_data[18]_INST_0_i_3_n_0 ),
        .I2(\read_data[23]_INST_0_i_6_n_0 ),
        .I3(addr[1]),
        .I4(\read_data[23]_INST_0_i_7_n_0 ),
        .I5(addr[0]),
        .O(\read_data[23]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000C3006AFF0000)) 
    \read_data[23]_INST_0_i_3 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[23]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \read_data[23]_INST_0_i_4 
       (.I0(addr[6]),
        .I1(addr[4]),
        .I2(addr[2]),
        .I3(addr[1]),
        .I4(addr[3]),
        .I5(addr[5]),
        .O(\read_data[23]_INST_0_i_4_n_0 ));
  MUXF7 \read_data[23]_INST_0_i_5 
       (.I0(\read_data[23]_INST_0_i_8_n_0 ),
        .I1(\read_data[23]_INST_0_i_9_n_0 ),
        .O(\read_data[23]_INST_0_i_5_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h0100100000802000)) 
    \read_data[23]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_9_n_0 ),
        .I2(\read_data[23]_INST_0_i_10_n_0 ),
        .I3(\read_data[23]_INST_0_i_11_n_0 ),
        .I4(\read_data[23]_INST_0_i_12_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[23]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000445444450)) 
    \read_data[23]_INST_0_i_7 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[23]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0001944500004444)) 
    \read_data[23]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(\read_data[20]_INST_0_i_7_n_0 ),
        .I2(\read_data[23]_INST_0_i_12_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[23]_INST_0_i_11_n_0 ),
        .I5(\read_data[20]_INST_0_i_9_n_0 ),
        .O(\read_data[23]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h020808080005CCC8)) 
    \read_data[23]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(\read_data[23]_INST_0_i_12_n_0 ),
        .I2(\read_data[23]_INST_0_i_11_n_0 ),
        .I3(\read_data[23]_INST_0_i_10_n_0 ),
        .I4(\read_data[20]_INST_0_i_9_n_0 ),
        .I5(\read_data[20]_INST_0_i_7_n_0 ),
        .O(\read_data[23]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[24]_INST_0 
       (.I0(\read_data[24]_INST_0_i_1_n_0 ),
        .I1(\read_data[31]_INST_0_i_2_n_0 ),
        .I2(\read_data[24]_INST_0_i_2_n_0 ),
        .I3(\read_data[31]_INST_0_i_4_n_0 ),
        .I4(\read_data[24]_INST_0_i_3_n_0 ),
        .O(read_data[24]));
  LUT6 #(
    .INIT(64'hE828E828EB2BE828)) 
    \read_data[24]_INST_0_i_1 
       (.I0(\read_data[24]_INST_0_i_4_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[24]_INST_0_i_5_n_0 ),
        .I4(\read_data[24]_INST_0_i_6_n_0 ),
        .I5(\read_data[31]_INST_0_i_8_n_0 ),
        .O(\read_data[24]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h6943C3C382800028)) 
    \read_data[24]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[24]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8141C3C3C3C3D7C3)) 
    \read_data[24]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[24]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000560001A800)) 
    \read_data[24]_INST_0_i_12 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[24]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hA9A8000001A85601)) 
    \read_data[24]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[24]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hA9A8000001A9A9A9)) 
    \read_data[24]_INST_0_i_14 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[24]_INST_0_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'h88800000)) 
    \read_data[24]_INST_0_i_15 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[3]),
        .O(\read_data[24]_INST_0_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'h1E)) 
    \read_data[24]_INST_0_i_16 
       (.I0(addr[1]),
        .I1(addr[0]),
        .I2(addr[2]),
        .O(\read_data[24]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[24]_INST_0_i_2 
       (.I0(\read_data[24]_INST_0_i_7_n_0 ),
        .I1(\read_data[24]_INST_0_i_8_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[24]_INST_0_i_9_n_0 ),
        .I5(\read_data[24]_INST_0_i_10_n_0 ),
        .O(\read_data[24]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0CA0F0A00CA000A0)) 
    \read_data[24]_INST_0_i_3 
       (.I0(\read_data[24]_INST_0_i_11_n_0 ),
        .I1(\read_data[24]_INST_0_i_12_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[24]_INST_0_i_13_n_0 ),
        .O(\read_data[24]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAEEEEAAA54444005)) 
    \read_data[24]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(\read_data[24]_INST_0_i_14_n_0 ),
        .I2(\read_data[24]_INST_0_i_15_n_0 ),
        .I3(addr[5]),
        .I4(addr[6]),
        .I5(\read_data[24]_INST_0_i_16_n_0 ),
        .O(\read_data[24]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0056565656000000)) 
    \read_data[24]_INST_0_i_5 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[24]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h1114333C333C333C)) 
    \read_data[24]_INST_0_i_6 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[24]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2800000000000028)) 
    \read_data[24]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[24]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h1110101444444444)) 
    \read_data[24]_INST_0_i_8 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[31]_INST_0_i_14_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[24]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h41438280402A402A)) 
    \read_data[24]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[24]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[25]_INST_0 
       (.I0(\read_data[25]_INST_0_i_1_n_0 ),
        .I1(\read_data[25]_INST_0_i_2_n_0 ),
        .I2(\read_data[31]_INST_0_i_2_n_0 ),
        .I3(\read_data[25]_INST_0_i_3_n_0 ),
        .I4(\read_data[31]_INST_0_i_4_n_0 ),
        .I5(\read_data[25]_INST_0_i_4_n_0 ),
        .O(read_data[25]));
  LUT5 #(
    .INIT(32'hEB2BE828)) 
    \read_data[25]_INST_0_i_1 
       (.I0(\read_data[25]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[25]_INST_0_i_6_n_0 ),
        .I4(\read_data[25]_INST_0_i_7_n_0 ),
        .O(\read_data[25]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h143C3C3C28284002)) 
    \read_data[25]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h2800414382800000)) 
    \read_data[25]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6943C3C38280402A)) 
    \read_data[25]_INST_0_i_12 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h015403FDFC03BC14)) 
    \read_data[25]_INST_0_i_13 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8014002800002815)) 
    \read_data[25]_INST_0_i_14 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hA800000000560001)) 
    \read_data[25]_INST_0_i_15 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[25]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFD0F0D0FF8000800)) 
    \read_data[25]_INST_0_i_2 
       (.I0(\read_data[31]_INST_0_i_8_n_0 ),
        .I1(\read_data[25]_INST_0_i_8_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[25]_INST_0_i_6_n_0 ),
        .I5(addr[2]),
        .O(\read_data[25]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[25]_INST_0_i_3 
       (.I0(\read_data[25]_INST_0_i_9_n_0 ),
        .I1(\read_data[25]_INST_0_i_10_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[25]_INST_0_i_11_n_0 ),
        .I5(\read_data[25]_INST_0_i_12_n_0 ),
        .O(\read_data[25]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0CA0FCA00CA00CA0)) 
    \read_data[25]_INST_0_i_4 
       (.I0(\read_data[25]_INST_0_i_13_n_0 ),
        .I1(\read_data[25]_INST_0_i_14_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[25]_INST_0_i_15_n_0 ),
        .O(\read_data[25]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000009FF99009)) 
    \read_data[25]_INST_0_i_5 
       (.I0(addr[1]),
        .I1(addr[2]),
        .I2(addr[6]),
        .I3(\read_data[31]_INST_0_i_6_n_0 ),
        .I4(\read_data[25]_INST_0_i_8_n_0 ),
        .I5(addr[0]),
        .O(\read_data[25]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5600000000565656)) 
    \read_data[25]_INST_0_i_6 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[25]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h3C3C3C3C3C3C7C3E)) 
    \read_data[25]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[25]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0808080000000080)) 
    \read_data[25]_INST_0_i_8 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[25]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0001010000000000)) 
    \read_data[25]_INST_0_i_9 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[31]_INST_0_i_14_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[25]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[26]_INST_0 
       (.I0(\read_data[26]_INST_0_i_1_n_0 ),
        .I1(\read_data[31]_INST_0_i_2_n_0 ),
        .I2(\read_data[26]_INST_0_i_2_n_0 ),
        .I3(\read_data[31]_INST_0_i_4_n_0 ),
        .I4(\read_data[26]_INST_0_i_3_n_0 ),
        .O(read_data[26]));
  LUT6 #(
    .INIT(64'hE3E3C0C3E0E0C0C3)) 
    \read_data[26]_INST_0_i_1 
       (.I0(\read_data[29]_INST_0_i_8_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[2]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[28]_INST_0_i_4_n_0 ),
        .O(\read_data[26]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[26]_INST_0_i_2 
       (.I0(\read_data[28]_INST_0_i_5_n_0 ),
        .I1(\read_data[26]_INST_0_i_4_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[26]_INST_0_i_5_n_0 ),
        .I5(\read_data[27]_INST_0_i_7_n_0 ),
        .O(\read_data[26]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFCA00CA0)) 
    \read_data[26]_INST_0_i_3 
       (.I0(\read_data[26]_INST_0_i_6_n_0 ),
        .I1(\read_data[26]_INST_0_i_7_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[26]_INST_0_i_8_n_0 ),
        .O(\read_data[26]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h02800000557FEA82)) 
    \read_data[26]_INST_0_i_4 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[26]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEBC3C3C3D7FFBFFD)) 
    \read_data[26]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[26]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000056AA5557AAA8)) 
    \read_data[26]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[26]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0014028028001400)) 
    \read_data[26]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[26]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFEA00004142416B)) 
    \read_data[26]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[26]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[27]_INST_0 
       (.I0(\read_data[27]_INST_0_i_1_n_0 ),
        .I1(\read_data[27]_INST_0_i_2_n_0 ),
        .I2(\read_data[31]_INST_0_i_2_n_0 ),
        .I3(\read_data[27]_INST_0_i_3_n_0 ),
        .I4(\read_data[31]_INST_0_i_4_n_0 ),
        .I5(\read_data[27]_INST_0_i_4_n_0 ),
        .O(read_data[27]));
  LUT5 #(
    .INIT(32'hEB2BE828)) 
    \read_data[27]_INST_0_i_1 
       (.I0(\read_data[27]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[29]_INST_0_i_7_n_0 ),
        .I4(\read_data[27]_INST_0_i_6_n_0 ),
        .O(\read_data[27]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0001FE0000000000)) 
    \read_data[27]_INST_0_i_10 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[27]_INST_0_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'h01010110)) 
    \read_data[27]_INST_0_i_11 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[2]),
        .I3(addr[1]),
        .I4(addr[0]),
        .O(\read_data[27]_INST_0_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'h57FFA800)) 
    \read_data[27]_INST_0_i_12 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .O(\read_data[27]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h9000900090000003)) 
    \read_data[27]_INST_0_i_13 
       (.I0(addr[4]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[1]),
        .I5(addr[0]),
        .O(\read_data[27]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \read_data[27]_INST_0_i_2 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .O(\read_data[27]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hEB2BE828)) 
    \read_data[27]_INST_0_i_3 
       (.I0(\read_data[27]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[29]_INST_0_i_7_n_0 ),
        .I4(\read_data[27]_INST_0_i_7_n_0 ),
        .O(\read_data[27]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0CA0F0A00CA000A0)) 
    \read_data[27]_INST_0_i_4 
       (.I0(\read_data[27]_INST_0_i_8_n_0 ),
        .I1(\read_data[27]_INST_0_i_9_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[27]_INST_0_i_10_n_0 ),
        .O(\read_data[27]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB08000000000B080)) 
    \read_data[27]_INST_0_i_5 
       (.I0(\read_data[27]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[27]_INST_0_i_12_n_0 ),
        .I3(\read_data[27]_INST_0_i_13_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[31]_INST_0_i_6_n_0 ),
        .O(\read_data[27]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hD7FFFFFFFFFFEBC3)) 
    \read_data[27]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[27]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h16BC3C3C7D7FEA82)) 
    \read_data[27]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[27]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0155A8005557AAA8)) 
    \read_data[27]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[27]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000005656000000)) 
    \read_data[27]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[27]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[28]_INST_0 
       (.I0(\read_data[28]_INST_0_i_1_n_0 ),
        .I1(\read_data[31]_INST_0_i_2_n_0 ),
        .I2(\read_data[28]_INST_0_i_2_n_0 ),
        .I3(\read_data[31]_INST_0_i_4_n_0 ),
        .I4(\read_data[28]_INST_0_i_3_n_0 ),
        .O(read_data[28]));
  LUT6 #(
    .INIT(64'h2323000320200003)) 
    \read_data[28]_INST_0_i_1 
       (.I0(\read_data[29]_INST_0_i_8_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[2]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[28]_INST_0_i_4_n_0 ),
        .O(\read_data[28]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0004040444545440)) 
    \read_data[28]_INST_0_i_10 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[31]_INST_0_i_14_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[28]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFEBFFFFFAAA9BEBD)) 
    \read_data[28]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[28]_INST_0_i_2 
       (.I0(\read_data[28]_INST_0_i_5_n_0 ),
        .I1(\read_data[29]_INST_0_i_12_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[28]_INST_0_i_6_n_0 ),
        .I5(\read_data[28]_INST_0_i_7_n_0 ),
        .O(\read_data[28]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[28]_INST_0_i_3 
       (.I0(\read_data[28]_INST_0_i_8_n_0 ),
        .I1(\read_data[28]_INST_0_i_9_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[28]_INST_0_i_10_n_0 ),
        .I5(\read_data[28]_INST_0_i_11_n_0 ),
        .O(\read_data[28]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEEBCCC3CCC3CCC3)) 
    \read_data[28]_INST_0_i_4 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[28]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4143C3C382800000)) 
    \read_data[28]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h143C3C3C28000000)) 
    \read_data[28]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h96BC3C3C7D7FFFD7)) 
    \read_data[28]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000001AAA80000)) 
    \read_data[28]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0015800028001400)) 
    \read_data[28]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[28]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[29]_INST_0 
       (.I0(\read_data[29]_INST_0_i_1_n_0 ),
        .I1(\read_data[29]_INST_0_i_2_n_0 ),
        .I2(\read_data[31]_INST_0_i_2_n_0 ),
        .I3(\read_data[29]_INST_0_i_3_n_0 ),
        .I4(\read_data[31]_INST_0_i_4_n_0 ),
        .I5(\read_data[29]_INST_0_i_4_n_0 ),
        .O(read_data[29]));
  LUT5 #(
    .INIT(32'hFCAF0CAF)) 
    \read_data[29]_INST_0_i_1 
       (.I0(\read_data[29]_INST_0_i_5_n_0 ),
        .I1(\read_data[29]_INST_0_i_6_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[29]_INST_0_i_7_n_0 ),
        .O(\read_data[29]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h294003C016BC6802)) 
    \read_data[29]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[29]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8014001580019401)) 
    \read_data[29]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[29]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000110000000)) 
    \read_data[29]_INST_0_i_12 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[31]_INST_0_i_14_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[29]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000444444440)) 
    \read_data[29]_INST_0_i_13 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[31]_INST_0_i_14_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[29]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h7EAA000055564142)) 
    \read_data[29]_INST_0_i_14 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[29]_INST_0_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \read_data[29]_INST_0_i_15 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .O(\read_data[29]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000F08888FFFF)) 
    \read_data[29]_INST_0_i_2 
       (.I0(\read_data[29]_INST_0_i_8_n_0 ),
        .I1(\read_data[31]_INST_0_i_8_n_0 ),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[0]),
        .I5(addr[1]),
        .O(\read_data[29]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF022FF00F022FF)) 
    \read_data[29]_INST_0_i_3 
       (.I0(\read_data[29]_INST_0_i_9_n_0 ),
        .I1(\read_data[31]_INST_0_i_8_n_0 ),
        .I2(\read_data[29]_INST_0_i_10_n_0 ),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(\read_data[29]_INST_0_i_7_n_0 ),
        .O(\read_data[29]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[29]_INST_0_i_4 
       (.I0(\read_data[29]_INST_0_i_11_n_0 ),
        .I1(\read_data[29]_INST_0_i_12_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[29]_INST_0_i_13_n_0 ),
        .I5(\read_data[29]_INST_0_i_14_n_0 ),
        .O(\read_data[29]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2A80000041438280)) 
    \read_data[29]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[29]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3D403FC03EBC3C00)) 
    \read_data[29]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[29]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h11155444)) 
    \read_data[29]_INST_0_i_7 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[29]_INST_0_i_15_n_0 ),
        .I4(addr[4]),
        .O(\read_data[29]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0808088080808080)) 
    \read_data[29]_INST_0_i_8 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[29]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0001A9A9A9A80000)) 
    \read_data[29]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[29]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFFBFB00000)) 
    \read_data[2]_INST_0 
       (.I0(\read_data[4]_INST_0_i_1_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[4]_INST_0_i_2_n_0 ),
        .I4(addr[8]),
        .I5(\read_data[2]_INST_0_i_1_n_0 ),
        .O(read_data[2]));
  MUXF8 \read_data[2]_INST_0_i_1 
       (.I0(\read_data[2]_INST_0_i_2_n_0 ),
        .I1(\read_data[2]_INST_0_i_3_n_0 ),
        .O(\read_data[2]_INST_0_i_1_n_0 ),
        .S(addr[7]));
  MUXF7 \read_data[2]_INST_0_i_2 
       (.I0(\read_data[2]_INST_0_i_4_n_0 ),
        .I1(\read_data[2]_INST_0_i_5_n_0 ),
        .O(\read_data[2]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[2]_INST_0_i_3 
       (.I0(\read_data[2]_INST_0_i_6_n_0 ),
        .I1(\read_data[2]_INST_0_i_7_n_0 ),
        .O(\read_data[2]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h2001191115D46000)) 
    \read_data[2]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAA00731)) 
    \read_data[2]_INST_0_i_5 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[3]),
        .I3(addr[4]),
        .I4(addr[6]),
        .I5(addr[0]),
        .O(\read_data[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0220966622006644)) 
    \read_data[2]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[5]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6DB7B796B795B795)) 
    \read_data[2]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[2]),
        .I3(addr[5]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[2]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[30]_INST_0 
       (.I0(\read_data[30]_INST_0_i_1_n_0 ),
        .I1(\read_data[30]_INST_0_i_2_n_0 ),
        .I2(\read_data[31]_INST_0_i_2_n_0 ),
        .I3(\read_data[30]_INST_0_i_3_n_0 ),
        .I4(\read_data[31]_INST_0_i_4_n_0 ),
        .I5(\read_data[30]_INST_0_i_4_n_0 ),
        .O(read_data[30]));
  LUT5 #(
    .INIT(32'hFCAF0CA0)) 
    \read_data[30]_INST_0_i_1 
       (.I0(\read_data[30]_INST_0_i_5_n_0 ),
        .I1(\read_data[30]_INST_0_i_6_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[30]_INST_0_i_7_n_0 ),
        .O(\read_data[30]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA801FFFE01A9A9A9)) 
    \read_data[30]_INST_0_i_10 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[30]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0014014180001400)) 
    \read_data[30]_INST_0_i_11 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[30]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000008080808000)) 
    \read_data[30]_INST_0_i_12 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[30]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h5657FFFFFFA9A800)) 
    \read_data[30]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[30]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0009090000)) 
    \read_data[30]_INST_0_i_2 
       (.I0(addr[4]),
        .I1(addr[3]),
        .I2(addr[2]),
        .I3(\read_data[30]_INST_0_i_8_n_0 ),
        .I4(addr[1]),
        .I5(addr[0]),
        .O(\read_data[30]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF022FF00F02200)) 
    \read_data[30]_INST_0_i_3 
       (.I0(\read_data[30]_INST_0_i_9_n_0 ),
        .I1(\read_data[31]_INST_0_i_8_n_0 ),
        .I2(\read_data[30]_INST_0_i_6_n_0 ),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(\read_data[30]_INST_0_i_7_n_0 ),
        .O(\read_data[30]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00F04400)) 
    \read_data[30]_INST_0_i_4 
       (.I0(\read_data[31]_INST_0_i_8_n_0 ),
        .I1(\read_data[30]_INST_0_i_10_n_0 ),
        .I2(\read_data[30]_INST_0_i_11_n_0 ),
        .I3(addr[1]),
        .I4(addr[0]),
        .O(\read_data[30]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hC003C003D403E803)) 
    \read_data[30]_INST_0_i_5 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[30]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2801828197C06AAA)) 
    \read_data[30]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[30]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBBF0F0BB88F0F088)) 
    \read_data[30]_INST_0_i_7 
       (.I0(\read_data[30]_INST_0_i_12_n_0 ),
        .I1(addr[0]),
        .I2(\read_data[24]_INST_0_i_6_n_0 ),
        .I3(\read_data[31]_INST_0_i_6_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[30]_INST_0_i_13_n_0 ),
        .O(\read_data[30]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEA83C003C003C003)) 
    \read_data[30]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[30]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0001FE01FE01A800)) 
    \read_data[30]_INST_0_i_9 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[30]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[31]_INST_0 
       (.I0(\read_data[31]_INST_0_i_1_n_0 ),
        .I1(\read_data[31]_INST_0_i_2_n_0 ),
        .I2(\read_data[31]_INST_0_i_3_n_0 ),
        .I3(\read_data[31]_INST_0_i_4_n_0 ),
        .I4(\read_data[31]_INST_0_i_5_n_0 ),
        .O(read_data[31]));
  LUT6 #(
    .INIT(64'h00009900007800FF)) 
    \read_data[31]_INST_0_i_1 
       (.I0(addr[3]),
        .I1(addr[4]),
        .I2(addr[5]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[31]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC0C0AFA0AFA0C0C0)) 
    \read_data[31]_INST_0_i_10 
       (.I0(\read_data[31]_INST_0_i_15_n_0 ),
        .I1(\read_data[31]_INST_0_i_16_n_0 ),
        .I2(addr[0]),
        .I3(\read_data[25]_INST_0_i_8_n_0 ),
        .I4(addr[6]),
        .I5(\read_data[31]_INST_0_i_6_n_0 ),
        .O(\read_data[31]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000001212121200)) 
    \read_data[31]_INST_0_i_11 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h01A8000000005600)) 
    \read_data[31]_INST_0_i_12 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[31]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0001FFFE000001A8)) 
    \read_data[31]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[31]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \read_data[31]_INST_0_i_14 
       (.I0(addr[0]),
        .I1(addr[1]),
        .O(\read_data[31]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCC14443CCC3CCC3)) 
    \read_data[31]_INST_0_i_15 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[1]),
        .I3(addr[0]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[31]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1818180404040484)) 
    \read_data[31]_INST_0_i_16 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(addr[2]),
        .O(\read_data[31]_INST_0_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \read_data[31]_INST_0_i_2 
       (.I0(addr[6]),
        .I1(\read_data[31]_INST_0_i_6_n_0 ),
        .I2(addr[7]),
        .I3(addr[8]),
        .O(\read_data[31]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF022FF00F02200)) 
    \read_data[31]_INST_0_i_3 
       (.I0(\read_data[31]_INST_0_i_7_n_0 ),
        .I1(\read_data[31]_INST_0_i_8_n_0 ),
        .I2(\read_data[31]_INST_0_i_9_n_0 ),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(\read_data[31]_INST_0_i_10_n_0 ),
        .O(\read_data[31]_INST_0_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \read_data[31]_INST_0_i_4 
       (.I0(\read_data[31]_INST_0_i_6_n_0 ),
        .I1(addr[6]),
        .I2(addr[7]),
        .O(\read_data[31]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00A0FC0000A00C00)) 
    \read_data[31]_INST_0_i_5 
       (.I0(\read_data[31]_INST_0_i_11_n_0 ),
        .I1(\read_data[31]_INST_0_i_12_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[31]_INST_0_i_8_n_0 ),
        .I5(\read_data[31]_INST_0_i_13_n_0 ),
        .O(\read_data[31]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8880000000000000)) 
    \read_data[31]_INST_0_i_6 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[31]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0001FFFE0001A800)) 
    \read_data[31]_INST_0_i_7 
       (.I0(addr[2]),
        .I1(addr[1]),
        .I2(addr[0]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[31]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \read_data[31]_INST_0_i_8 
       (.I0(\read_data[31]_INST_0_i_6_n_0 ),
        .I1(addr[6]),
        .O(\read_data[31]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4143828015558000)) 
    \read_data[31]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[31]_INST_0_i_14_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[31]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[3]_INST_0 
       (.I0(\read_data[3]_INST_0_i_1_n_0 ),
        .I1(\read_data[3]_INST_0_i_2_n_0 ),
        .O(read_data[3]),
        .S(addr[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[3]_INST_0_i_1 
       (.I0(\read_data[3]_INST_0_i_3_n_0 ),
        .I1(\read_data[3]_INST_0_i_4_n_0 ),
        .I2(addr[7]),
        .I3(\read_data[3]_INST_0_i_5_n_0 ),
        .I4(addr[1]),
        .I5(\read_data[3]_INST_0_i_6_n_0 ),
        .O(\read_data[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFA0A0C0C0C0C0)) 
    \read_data[3]_INST_0_i_2 
       (.I0(\read_data[3]_INST_0_i_7_n_0 ),
        .I1(\read_data[3]_INST_0_i_4_n_0 ),
        .I2(addr[7]),
        .I3(addr[2]),
        .I4(addr[0]),
        .I5(addr[1]),
        .O(\read_data[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h488888888FF0F7F0)) 
    \read_data[3]_INST_0_i_3 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[5]),
        .I3(addr[4]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000408)) 
    \read_data[3]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(addr[4]),
        .I2(addr[5]),
        .I3(addr[2]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000040)) 
    \read_data[3]_INST_0_i_5 
       (.I0(addr[6]),
        .I1(addr[4]),
        .I2(addr[5]),
        .I3(addr[2]),
        .I4(addr[3]),
        .I5(addr[0]),
        .O(\read_data[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00011D55D1100000)) 
    \read_data[3]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4CCCCCCCCFF4F7F4)) 
    \read_data[3]_INST_0_i_7 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[5]),
        .I3(addr[4]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8F80FFFF8F800000)) 
    \read_data[4]_INST_0 
       (.I0(\read_data[4]_INST_0_i_1_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[4]_INST_0_i_2_n_0 ),
        .I4(addr[8]),
        .I5(\read_data[4]_INST_0_i_3_n_0 ),
        .O(read_data[4]));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'h8000FFFF)) 
    \read_data[4]_INST_0_i_1 
       (.I0(addr[5]),
        .I1(addr[3]),
        .I2(addr[4]),
        .I3(addr[6]),
        .I4(addr[2]),
        .O(\read_data[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \read_data[4]_INST_0_i_2 
       (.I0(addr[6]),
        .I1(addr[3]),
        .I2(addr[5]),
        .I3(addr[4]),
        .I4(addr[0]),
        .O(\read_data[4]_INST_0_i_2_n_0 ));
  MUXF8 \read_data[4]_INST_0_i_3 
       (.I0(\read_data[4]_INST_0_i_4_n_0 ),
        .I1(\read_data[4]_INST_0_i_5_n_0 ),
        .O(\read_data[4]_INST_0_i_3_n_0 ),
        .S(addr[7]));
  MUXF7 \read_data[4]_INST_0_i_4 
       (.I0(\read_data[4]_INST_0_i_6_n_0 ),
        .I1(\read_data[4]_INST_0_i_7_n_0 ),
        .O(\read_data[4]_INST_0_i_4_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[4]_INST_0_i_5 
       (.I0(\read_data[4]_INST_0_i_8_n_0 ),
        .I1(\read_data[4]_INST_0_i_9_n_0 ),
        .O(\read_data[4]_INST_0_i_5_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h3010100002008084)) 
    \read_data[4]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[5]),
        .I3(addr[2]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA2AAAAE4746A)) 
    \read_data[4]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(addr[5]),
        .I2(addr[2]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[6]),
        .O(\read_data[4]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000144600004444)) 
    \read_data[4]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[5]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h3E82EC22EE22EE22)) 
    \read_data[4]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[4]),
        .O(\read_data[4]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[5]_INST_0 
       (.I0(\read_data[5]_INST_0_i_1_n_0 ),
        .I1(\read_data[5]_INST_0_i_2_n_0 ),
        .O(read_data[5]),
        .S(addr[8]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \read_data[5]_INST_0_i_1 
       (.I0(\read_data[5]_INST_0_i_3_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[5]_INST_0_i_4_n_0 ),
        .I4(addr[7]),
        .I5(\read_data[5]_INST_0_i_5_n_0 ),
        .O(\read_data[5]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFA0CFCFFFA0C0C0)) 
    \read_data[5]_INST_0_i_2 
       (.I0(\read_data[5]_INST_0_i_3_n_0 ),
        .I1(\read_data[5]_INST_0_i_6_n_0 ),
        .I2(addr[7]),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(\read_data[5]_INST_0_i_7_n_0 ),
        .O(\read_data[5]_INST_0_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'h006E)) 
    \read_data[5]_INST_0_i_3 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[6]),
        .O(\read_data[5]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8222000029909290)) 
    \read_data[5]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(addr[2]),
        .I2(addr[5]),
        .I3(addr[4]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[5]_INST_0_i_4_n_0 ));
  MUXF7 \read_data[5]_INST_0_i_5 
       (.I0(\read_data[5]_INST_0_i_8_n_0 ),
        .I1(\read_data[5]_INST_0_i_9_n_0 ),
        .O(\read_data[5]_INST_0_i_5_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'hE2A2A0A061919080)) 
    \read_data[5]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[4]),
        .I4(addr[5]),
        .I5(addr[2]),
        .O(\read_data[5]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB888000088880000)) 
    \read_data[5]_INST_0_i_7 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[4]),
        .I3(addr[5]),
        .I4(addr[3]),
        .I5(addr[6]),
        .O(\read_data[5]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200411045)) 
    \read_data[5]_INST_0_i_8 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[2]),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[4]),
        .O(\read_data[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88888000000ECEC0)) 
    \read_data[5]_INST_0_i_9 
       (.I0(addr[0]),
        .I1(addr[5]),
        .I2(addr[2]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[6]),
        .O(\read_data[5]_INST_0_i_9_n_0 ));
  MUXF7 \read_data[6]_INST_0 
       (.I0(\read_data[6]_INST_0_i_1_n_0 ),
        .I1(\read_data[6]_INST_0_i_2_n_0 ),
        .O(read_data[6]),
        .S(addr[8]));
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data[6]_INST_0_i_1 
       (.I0(\read_data[6]_INST_0_i_3_n_0 ),
        .I1(\read_data[6]_INST_0_i_4_n_0 ),
        .I2(addr[7]),
        .I3(\read_data[6]_INST_0_i_5_n_0 ),
        .I4(addr[1]),
        .O(\read_data[6]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data[6]_INST_0_i_2 
       (.I0(\read_data[6]_INST_0_i_3_n_0 ),
        .I1(\read_data[6]_INST_0_i_6_n_0 ),
        .I2(addr[7]),
        .I3(\read_data[6]_INST_0_i_7_n_0 ),
        .I4(addr[1]),
        .O(\read_data[6]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3E02EC22EE22CC00)) 
    \read_data[6]_INST_0_i_3 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[4]),
        .O(\read_data[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h820000222E1BE010)) 
    \read_data[6]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(addr[2]),
        .I2(addr[5]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[6]),
        .O(\read_data[6]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0002002226201066)) 
    \read_data[6]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[4]),
        .O(\read_data[6]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8330002022A05D7D)) 
    \read_data[6]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[4]),
        .I3(addr[5]),
        .I4(addr[3]),
        .I5(addr[2]),
        .O(\read_data[6]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE0A040000A0A5555)) 
    \read_data[6]_INST_0_i_7 
       (.I0(addr[0]),
        .I1(addr[5]),
        .I2(addr[4]),
        .I3(addr[6]),
        .I4(addr[2]),
        .I5(addr[3]),
        .O(\read_data[6]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[7]_INST_0 
       (.I0(\read_data[7]_INST_0_i_1_n_0 ),
        .I1(addr[8]),
        .I2(\read_data[7]_INST_0_i_2_n_0 ),
        .I3(addr[7]),
        .I4(\read_data[7]_INST_0_i_3_n_0 ),
        .O(read_data[7]));
  LUT6 #(
    .INIT(64'h1400AA005000AA55)) 
    \read_data[7]_INST_0_i_1 
       (.I0(addr[1]),
        .I1(addr[3]),
        .I2(addr[5]),
        .I3(addr[0]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[7]_INST_0_i_1_n_0 ));
  MUXF7 \read_data[7]_INST_0_i_2 
       (.I0(\read_data[7]_INST_0_i_4_n_0 ),
        .I1(\read_data[7]_INST_0_i_5_n_0 ),
        .O(\read_data[7]_INST_0_i_2_n_0 ),
        .S(addr[1]));
  MUXF7 \read_data[7]_INST_0_i_3 
       (.I0(\read_data[7]_INST_0_i_6_n_0 ),
        .I1(\read_data[7]_INST_0_i_7_n_0 ),
        .O(\read_data[7]_INST_0_i_3_n_0 ),
        .S(addr[1]));
  LUT6 #(
    .INIT(64'h020808080005CCC8)) 
    \read_data[7]_INST_0_i_4 
       (.I0(addr[0]),
        .I1(addr[5]),
        .I2(addr[2]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[6]),
        .O(\read_data[7]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0001944500004444)) 
    \read_data[7]_INST_0_i_5 
       (.I0(addr[0]),
        .I1(addr[6]),
        .I2(addr[5]),
        .I3(addr[3]),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[7]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0100100000802000)) 
    \read_data[7]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[7]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011140010)) 
    \read_data[7]_INST_0_i_7 
       (.I0(addr[6]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[2]),
        .I4(addr[5]),
        .I5(addr[0]),
        .O(\read_data[7]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \read_data[8]_INST_0 
       (.I0(\read_data[8]_INST_0_i_1_n_0 ),
        .I1(\read_data[15]_INST_0_i_2_n_0 ),
        .I2(\read_data[8]_INST_0_i_2_n_0 ),
        .I3(\read_data[15]_INST_0_i_4_n_0 ),
        .I4(\read_data[8]_INST_0_i_3_n_0 ),
        .O(read_data[8]));
  LUT6 #(
    .INIT(64'hFF0CAAFF000CAA00)) 
    \read_data[8]_INST_0_i_1 
       (.I0(\read_data[8]_INST_0_i_4_n_0 ),
        .I1(\read_data[8]_INST_0_i_5_n_0 ),
        .I2(\read_data[15]_INST_0_i_9_n_0 ),
        .I3(addr[0]),
        .I4(addr[1]),
        .I5(\read_data[8]_INST_0_i_6_n_0 ),
        .O(\read_data[8]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1110101444444444)) 
    \read_data[8]_INST_0_i_10 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[15]_INST_0_i_16_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[8]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h9580000015806A15)) 
    \read_data[8]_INST_0_i_11 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[8]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8141C3C3C3C3D7C3)) 
    \read_data[8]_INST_0_i_12 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[8]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000006A00158000)) 
    \read_data[8]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h9580000015959595)) 
    \read_data[8]_INST_0_i_14 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[8]_INST_0_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \read_data[8]_INST_0_i_15 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(addr[3]),
        .O(\read_data[8]_INST_0_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \read_data[8]_INST_0_i_16 
       (.I0(addr[0]),
        .I1(addr[1]),
        .I2(addr[2]),
        .O(\read_data[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[8]_INST_0_i_2 
       (.I0(\read_data[8]_INST_0_i_7_n_0 ),
        .I1(\read_data[8]_INST_0_i_8_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[8]_INST_0_i_9_n_0 ),
        .I5(\read_data[8]_INST_0_i_10_n_0 ),
        .O(\read_data[8]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC303C000C808C808)) 
    \read_data[8]_INST_0_i_3 
       (.I0(\read_data[8]_INST_0_i_11_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(\read_data[8]_INST_0_i_12_n_0 ),
        .I4(\read_data[8]_INST_0_i_13_n_0 ),
        .I5(\read_data[15]_INST_0_i_9_n_0 ),
        .O(\read_data[8]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h006A6A6A6A000000)) 
    \read_data[8]_INST_0_i_4 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[8]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h14443CCC3CCC3CCC)) 
    \read_data[8]_INST_0_i_5 
       (.I0(addr[5]),
        .I1(addr[2]),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(addr[3]),
        .I5(addr[4]),
        .O(\read_data[8]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAEEEEAAA54444005)) 
    \read_data[8]_INST_0_i_6 
       (.I0(addr[0]),
        .I1(\read_data[8]_INST_0_i_14_n_0 ),
        .I2(\read_data[8]_INST_0_i_15_n_0 ),
        .I3(addr[5]),
        .I4(addr[6]),
        .I5(\read_data[8]_INST_0_i_16_n_0 ),
        .O(\read_data[8]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h41438280402A402A)) 
    \read_data[8]_INST_0_i_7 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[8]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h6943C3C382800028)) 
    \read_data[8]_INST_0_i_8 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2800000000000028)) 
    \read_data[8]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[8]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data[9]_INST_0 
       (.I0(\read_data[9]_INST_0_i_1_n_0 ),
        .I1(\read_data[9]_INST_0_i_2_n_0 ),
        .I2(\read_data[15]_INST_0_i_2_n_0 ),
        .I3(\read_data[9]_INST_0_i_3_n_0 ),
        .I4(\read_data[15]_INST_0_i_4_n_0 ),
        .I5(\read_data[9]_INST_0_i_4_n_0 ),
        .O(read_data[9]));
  LUT5 #(
    .INIT(32'hFCAF0CA0)) 
    \read_data[9]_INST_0_i_1 
       (.I0(\read_data[9]_INST_0_i_5_n_0 ),
        .I1(\read_data[9]_INST_0_i_6_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[9]_INST_0_i_7_n_0 ),
        .O(\read_data[9]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h6943C3C38280402A)) 
    \read_data[9]_INST_0_i_10 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0001010000000000)) 
    \read_data[9]_INST_0_i_11 
       (.I0(addr[6]),
        .I1(addr[5]),
        .I2(addr[3]),
        .I3(\read_data[15]_INST_0_i_16_n_0 ),
        .I4(addr[2]),
        .I5(addr[4]),
        .O(\read_data[9]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h143C3C3C28284002)) 
    \read_data[9]_INST_0_i_12 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h80000000006A0015)) 
    \read_data[9]_INST_0_i_13 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[9]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h015403FDFC03BC14)) 
    \read_data[9]_INST_0_i_14 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8014002800002815)) 
    \read_data[9]_INST_0_i_15 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3B0B380B3808380B)) 
    \read_data[9]_INST_0_i_2 
       (.I0(\read_data[9]_INST_0_i_5_n_0 ),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[2]),
        .I4(\read_data[15]_INST_0_i_9_n_0 ),
        .I5(\read_data[9]_INST_0_i_8_n_0 ),
        .O(\read_data[9]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFCAF0CAFFCA00CA0)) 
    \read_data[9]_INST_0_i_3 
       (.I0(\read_data[9]_INST_0_i_9_n_0 ),
        .I1(\read_data[9]_INST_0_i_10_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[9]_INST_0_i_11_n_0 ),
        .I5(\read_data[9]_INST_0_i_12_n_0 ),
        .O(\read_data[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF04F004FF0400040)) 
    \read_data[9]_INST_0_i_4 
       (.I0(\read_data[15]_INST_0_i_9_n_0 ),
        .I1(\read_data[9]_INST_0_i_13_n_0 ),
        .I2(addr[0]),
        .I3(addr[1]),
        .I4(\read_data[9]_INST_0_i_14_n_0 ),
        .I5(\read_data[9]_INST_0_i_15_n_0 ),
        .O(\read_data[9]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6A000000006A6A6A)) 
    \read_data[9]_INST_0_i_5 
       (.I0(addr[2]),
        .I1(addr[0]),
        .I2(addr[1]),
        .I3(addr[3]),
        .I4(addr[4]),
        .I5(addr[5]),
        .O(\read_data[9]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3C3C3C3C3C3C7C3E)) 
    \read_data[9]_INST_0_i_6 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT5 #(
    .INIT(32'h00007D41)) 
    \read_data[9]_INST_0_i_7 
       (.I0(addr[2]),
        .I1(addr[6]),
        .I2(\read_data[15]_INST_0_i_6_n_0 ),
        .I3(\read_data[9]_INST_0_i_8_n_0 ),
        .I4(addr[0]),
        .O(\read_data[9]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000808080)) 
    \read_data[9]_INST_0_i_8 
       (.I0(addr[5]),
        .I1(addr[4]),
        .I2(addr[3]),
        .I3(addr[1]),
        .I4(addr[0]),
        .I5(addr[2]),
        .O(\read_data[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2800414382800000)) 
    \read_data[9]_INST_0_i_9 
       (.I0(addr[4]),
        .I1(addr[2]),
        .I2(\read_data[15]_INST_0_i_16_n_0 ),
        .I3(addr[3]),
        .I4(addr[5]),
        .I5(addr[6]),
        .O(\read_data[9]_INST_0_i_9_n_0 ));
endmodule
